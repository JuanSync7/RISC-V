//=============================================================================
// Company: Sondrel Ltd
// Author: DesignAI (designai@sondrel.com)
// Created: 2025-01-27
//
// File: tilelink_adapter.sv
// Module: tilelink_adapter
//
// Project Name: RISC-V RV32IM Core
// Target Devices: ASIC/FPGA
// Tool Versions: VCS 2020.03, ModelSim 2021.1
// Verification Status: Not Verified
// Quality Status: Draft
//
// Description:
//   TileLink protocol adapter that translates between the generic memory
//   interface and TileLink protocol. Supports TileLink Uncached (TL-UL)
//   and TileLink Cached (TL-C) protocols for RISC-V ecosystem integration.
//   Updated to use proper interface.
//=============================================================================

`timescale 1ns/1ps
`default_nettype none

// AI_TAG: FEATURE - TileLink protocol translation from generic memory interface using proper interface
// AI_TAG: FEATURE - Support for TL-UL (Uncached) and TL-C (Cached) operations
// AI_TAG: FEATURE - Transaction ID tracking and response matching
// AI_TAG: FEATURE - Burst support for cache line operations using TileLink interface

import riscv_config_pkg::*;
import riscv_types_pkg::*;
import riscv_protocol_types_pkg::*;
import riscv_core_pkg::*;

module tilelink_adapter #(
    parameter integer ADDR_WIDTH = 32,         // AI_TAG: PARAM_DESC - Address bus width
                                               // AI_TAG: PARAM_USAGE - Must match tilelink_if parameter
                                               // AI_TAG: PARAM_CONSTRAINTS - Must match tilelink_if parameter
    parameter integer DATA_WIDTH = 32,         // AI_TAG: PARAM_DESC - Data bus width
                                               // AI_TAG: PARAM_USAGE - Must match tilelink_if parameter
                                               // AI_TAG: PARAM_CONSTRAINTS - Must match tilelink_if parameter
    parameter integer SOURCE_WIDTH = 8,        // AI_TAG: PARAM_DESC - TileLink source ID width
                                               // AI_TAG: PARAM_USAGE - Must match tilelink_if parameter
                                               // AI_TAG: PARAM_CONSTRAINTS - Must match tilelink_if parameter
    parameter integer SINK_WIDTH = 8,          // AI_TAG: PARAM_DESC - TileLink sink ID width
                                               // AI_TAG: PARAM_USAGE - Must match tilelink_if parameter
                                               // AI_TAG: PARAM_CONSTRAINTS - Must match tilelink_if parameter
    parameter integer SIZE_WIDTH = 3,          // AI_TAG: PARAM_DESC - TileLink size width
                                               // AI_TAG: PARAM_USAGE - Must match tilelink_if parameter
                                               // AI_TAG: PARAM_CONSTRAINTS - Must match tilelink_if parameter
    parameter integer MAX_OUTSTANDING = 16     // AI_TAG: PARAM_DESC - Maximum outstanding transactions
                                               // AI_TAG: PARAM_USAGE - Sets transaction table size
                                               // AI_TAG: PARAM_CONSTRAINTS - Must be power of 2, max 256
) (
    input  logic        clk_i,     // AI_TAG: PORT_DESC - System clock
                                   // AI_TAG: PORT_CLK_DOMAIN - clk_i
    input  logic        rst_ni,    // AI_TAG: PORT_DESC - Asynchronous active-low reset
                                   // AI_TAG: PORT_CLK_DOMAIN - clk_i (async assert)
                                   // AI_TAG: PORT_TIMING - Asynchronous

    // Generic memory interface
    // AI_TAG: IF_TYPE - Generic Memory Interface (slave)
    // AI_TAG: IF_DESC - Protocol-agnostic memory interface
    // AI_TAG: IF_CLOCKING - clk_i
    // AI_TAG: IF_RESET - rst_ni
    memory_req_rsp_if.slave mem_if,

    // TileLink Interface - Using proper interface
    // AI_TAG: IF_TYPE - TileLink Manager (Client)
    // AI_TAG: IF_MODPORT - manager
    // AI_TAG: IF_PROTOCOL_VERSION - TileLink Uncached (TL-UL)
    // AI_TAG: IF_DESC - TileLink interface for open-source ecosystem compatibility
    // AI_TAG: IF_DATA_WIDTHS - Data: parameterized, Addr: parameterized, Source: parameterized
    // AI_TAG: IF_CLOCKING - clk_i via tl_if.clk connection
    // AI_TAG: IF_RESET - rst_ni via tl_if.reset_n connection
    tilelink_if.manager tl_if
);

    // AI_TAG: INTERNAL_BLOCK - TransactionTracker - Manages outstanding TileLink transactions
    // AI_TAG: INTERNAL_BLOCK - StateMachine - Controls TileLink transaction flow
    // AI_TAG: INTERNAL_BLOCK - ProtocolConverter - Converts between memory and TileLink protocols

    // Connect interface clock and reset
    assign tl_if.clk = clk_i;
    assign tl_if.reset_n = rst_ni;

    // AI_TAG: DATAPATH_DESC - Memory requests are converted to TileLink A-channel requests, D-channel responses are converted back

    // Import protocol constants package for TileLink opcodes
    import riscv_protocol_constants_pkg::*;
    import riscv_qos_pkg::*;

    //-----
    // Transaction Tracking
    //-----
    // AI_TAG: INTERNAL_STORAGE - Transaction table for tracking outstanding requests
    // AI_TAG: INTERNAL_STORAGE_TYPE - Transaction table - Memory array
    // AI_TAG: INTERNAL_STORAGE_ACCESS - Transaction table - FSM controlled
    typedef struct packed {
        logic                       valid;
        logic                       is_write;
        logic [ADDR_WIDTH-1:0]      addr;
        logic [DATA_WIDTH-1:0]      data;
        logic [(DATA_WIDTH/8)-1:0]  mask;
        logic [15:0]                mem_req_id;  // Original memory request ID
        logic                       response_pending;
        logic [SOURCE_WIDTH-1:0]    tl_source_id;
    } transaction_entry_t;

    transaction_entry_t transaction_table [MAX_OUTSTANDING-1:0];
    logic [SOURCE_WIDTH-1:0] next_source_id;
    logic [SOURCE_WIDTH-1:0] allocated_source_id;
    logic                    txn_alloc_valid;

    // AI_TAG: FSM_NAME - tilelink_adapter_fsm
    // AI_TAG: FSM_PURPOSE - tilelink_adapter_fsm - Controls TileLink transaction flow and state management
    // AI_TAG: FSM_ENCODING - tilelink_adapter_fsm - binary
    // AI_TAG: FSM_RESET_STATE - tilelink_adapter_fsm - IDLE
    typedef enum logic [2:0] {
        IDLE,               // AI_TAG: FSM_STATE - IDLE - Waiting for request or checking responses
        SEND_REQUEST,       // AI_TAG: FSM_STATE - SEND_REQUEST - Sending TileLink A-channel request
        WAIT_RESPONSE,      // AI_TAG: FSM_STATE - WAIT_RESPONSE - Waiting for TileLink D-channel response
        SEND_GENERIC_RSP    // AI_TAG: FSM_STATE - SEND_GENERIC_RSP - Sending response to memory interface
    } state_e;

    state_e current_state_q, next_state_c;

    //-----
    // Internal Signals
    //-----
    logic can_accept_request;
    logic [SOURCE_WIDTH-1:0] free_source_id;
    logic found_free_slot;
    logic [SIZE_WIDTH-1:0] transfer_size;
    logic [SOURCE_WIDTH-1:0] completed_source_id;
    logic completed_txn_valid;

    //-----
    // Transfer size calculation
    //-----
    always_comb begin : proc_transfer_size
        // Calculate log2 of transfer size in bytes based on memory request size
        case (mem_if.req.size)
            3'd0: transfer_size = 3'd0; // 1 byte
            3'd1: transfer_size = 3'd1; // 2 bytes
            3'd2: transfer_size = 3'd2; // 4 bytes
            3'd3: transfer_size = 3'd3; // 8 bytes
            default: transfer_size = 3'd2; // Default to 4 bytes
        endcase
    end

    //-----
    // Source ID Management
    //-----
    always_ff @(posedge clk_i or negedge rst_ni) begin : proc_source_id_counter
        if (!rst_ni) begin
            next_source_id <= '0;
        end else if (txn_alloc_valid) begin
            next_source_id <= next_source_id + 1;
        end
    end

    // Find free transaction slot
    always_comb begin : proc_find_free_slot
        found_free_slot = 1'b0;
        free_source_id = '0;
        
        for (int i = 0; i < MAX_OUTSTANDING; i++) begin
            if (!transaction_table[i].valid) begin
                found_free_slot = 1'b1;
                free_source_id = i[SOURCE_WIDTH-1:0];
                break;
            end
        end
    end

    // Find completed transaction for response
    always_comb begin : proc_find_completed_txn
        completed_txn_valid = 1'b0;
        completed_source_id = '0;
        
        for (int i = 0; i < MAX_OUTSTANDING; i++) begin
            if (transaction_table[i].valid && !transaction_table[i].response_pending) begin
                completed_txn_valid = 1'b1;
                completed_source_id = i[SOURCE_WIDTH-1:0];
                break;
            end
        end
    end

    assign can_accept_request = found_free_slot;
    assign allocated_source_id = free_source_id;

    // AI_TAG: FSM_TRANSITION - tilelink_adapter_fsm: IDLE -> SEND_REQUEST when (mem_if.req_valid && can_accept_request)
    // AI_TAG: FSM_TRANSITION - tilelink_adapter_fsm: SEND_REQUEST -> WAIT_RESPONSE when (tl_if.a_valid && tl_if.a_ready)
    // AI_TAG: FSM_TRANSITION - tilelink_adapter_fsm: WAIT_RESPONSE -> IDLE when response processed
    // AI_TAG: FSM_TRANSITION - tilelink_adapter_fsm: SEND_GENERIC_RSP -> IDLE when (mem_if.rsp_ready)

    //-----
    // Main FSM
    //-----
    always_ff @(posedge clk_i or negedge rst_ni) begin : proc_fsm_state
        if (!rst_ni) begin
            current_state_q <= IDLE;
            for (int i = 0; i < MAX_OUTSTANDING; i++) begin
                transaction_table[i] <= '0;
            end
        end else begin
            current_state_q <= next_state_c;
            
            // Handle transaction allocation
            if (txn_alloc_valid) begin
                transaction_table[allocated_source_id].valid <= 1'b1;
                transaction_table[allocated_source_id].is_write <= mem_if.req.write;
                transaction_table[allocated_source_id].addr <= mem_if.req.addr;
                transaction_table[allocated_source_id].data <= mem_if.req.data;
                transaction_table[allocated_source_id].mask <= mem_if.req.strb[(DATA_WIDTH/8)-1:0];
                transaction_table[allocated_source_id].mem_req_id <= mem_if.req.id;
                transaction_table[allocated_source_id].response_pending <= 1'b1;
                transaction_table[allocated_source_id].tl_source_id <= next_source_id;
            end
            
            // Handle response reception
            if (tl_if.d_valid && tl_if.d_ready) begin
                for (int i = 0; i < MAX_OUTSTANDING; i++) begin
                    if (transaction_table[i].valid && 
                        transaction_table[i].tl_source_id == tl_if.d_source) begin
                        transaction_table[i].response_pending <= 1'b0;
                        break;
                    end
                end
            end
            
            // Clear completed transactions
            if (mem_if.rsp_valid && mem_if.rsp_ready) begin
                transaction_table[completed_source_id].valid <= 1'b0;
            end
        end
    end

    always_comb begin : proc_fsm_logic
        next_state_c = current_state_q;
        
        // Default memory interface outputs
        mem_if.req_ready = 1'b0;
        mem_if.rsp_valid = 1'b0;
        mem_if.rsp = '0;
        
        // Default TileLink interface outputs
        tl_if.a_valid = 1'b0;
        tl_if.a_opcode = '0;
        tl_if.a_param = '0;
        tl_if.a_size = transfer_size;
        tl_if.a_source = '0;
        tl_if.a_address = '0;
        tl_if.a_mask = '0;
        tl_if.a_data = '0;
        tl_if.a_corrupt = 1'b0;
        tl_if.a_user = '0;
        
        tl_if.d_ready = 1'b1;  // Always ready to accept responses
        
        txn_alloc_valid = 1'b0;

        case (current_state_q)
            IDLE: begin
                mem_if.req_ready = can_accept_request;
                
                if (mem_if.req_valid && can_accept_request) begin
                    txn_alloc_valid = 1'b1;
                    next_state_c = SEND_REQUEST;
                end else if (completed_txn_valid) begin
                    next_state_c = SEND_GENERIC_RSP;
                end
            end

            SEND_REQUEST: begin
                tl_if.a_valid = 1'b1;
                tl_if.a_source = next_source_id;
                tl_if.a_address = mem_if.req.addr;
                tl_if.a_size = transfer_size;
                tl_if.a_mask = mem_if.req.strb[(DATA_WIDTH/8)-1:0];
                
                if (mem_if.req.write) begin
                    // Determine if full or partial write based on strobe pattern
                    if (mem_if.req.strb == {(DATA_WIDTH/8){1'b1}}) begin
                        tl_if.a_opcode = TL_A_PutFullData;
                    end else begin
                        tl_if.a_opcode = TL_A_PutPartialData;
                    end
                    tl_if.a_data = mem_if.req.data;
                end else begin
                    tl_if.a_opcode = TL_A_Get;
                    tl_if.a_data = RESET_VALUE_32BIT;
                end
                
                // Set default parameters
                tl_if.a_param = TL_PARAM_NO_PARAM;  // No specific parameters for TL-UL
                
                // QoS Assignment Logic - TileLink priority mapping
                logic [3:0] dynamic_qos_level;
                qos_transaction_type_e transaction_type;
                
                // Determine transaction type based on address and access pattern
                if (mem_if.req.addr >= 32'h0000_0000 && mem_if.req.addr < 32'h0000_1000) begin
                    transaction_type = QOS_TYPE_EXCEPTION;  // Exception vectors
                end else if (!mem_if.req.write && (mem_if.req.addr[1:0] == 2'b00)) begin
                    transaction_type = QOS_TYPE_INSTR_FETCH; // Likely instruction fetch
                end else if (mem_if.req.write || mem_if.req.strb != 4'hF) begin
                    transaction_type = QOS_TYPE_DATA_ACCESS; // Data access
                end else if (mem_if.req.addr >= 32'hF000_0000) begin
                    transaction_type = QOS_TYPE_PERIPHERAL;  // Peripheral space
                end else begin
                    transaction_type = QOS_TYPE_CACHE_FILL;  // Default to cache fill
                end
                
                // Dynamic QoS level assignment (embedded in user field for TileLink)
                dynamic_qos_level = get_qos_level(transaction_type);
                tl_if.a_user[3:0] = dynamic_qos_level;   // QoS in user field
                tl_if.a_user[7:4] = 4'h0; // Reserved user bits
                
                if (tl_if.a_ready) begin
                    next_state_c = WAIT_RESPONSE;
                end
            end

            WAIT_RESPONSE: begin
                // Wait for response, handled by transaction table updates
                if (completed_txn_valid) begin
                    next_state_c = SEND_GENERIC_RSP;
                end else begin
                    next_state_c = IDLE;
                end
            end

            SEND_GENERIC_RSP: begin
                mem_if.rsp_valid = 1'b1;
                mem_if.rsp.id = transaction_table[completed_source_id].mem_req_id;
                mem_if.rsp.last = 1'b1;
                
                if (!transaction_table[completed_source_id].is_write) begin
                    // Read response - get data from TileLink D-channel
                    if (tl_if.d_valid && 
                        tl_if.d_source == transaction_table[completed_source_id].tl_source_id) begin
                        mem_if.rsp.data = tl_if.d_data;
                        mem_if.rsp.error = tl_if.d_denied || tl_if.d_corrupt;
                    end else begin
                        mem_if.rsp.data = '0;
                        mem_if.rsp.error = 1'b0;
                    end
                end else begin
                    // Write response - no data needed
                    mem_if.rsp.data = '0;
                    mem_if.rsp.error = tl_if.d_denied || tl_if.d_corrupt;
                end
                
                if (mem_if.rsp_ready) begin
                    next_state_c = IDLE;
                end
            end

            default: begin
                next_state_c = IDLE;
            end
        endcase
    end

    //-----
    // TileLink Response Validation
    //-----
    logic valid_response_opcode;
    
    always_comb begin : proc_response_validation
        valid_response_opcode = 1'b0;
        case (tl_if.d_opcode)
            TL_AccessAck, TL_AccessAckData: valid_response_opcode = 1'b1;
            default: valid_response_opcode = 1'b0;
        endcase
    end

    // AI_TAG: ASSERTION - a_transaction_table_no_overflow: Transaction table should not overflow
    // AI_TAG: ASSERTION_TYPE - Simulation
    // AI_TAG: ASSERTION_SEVERITY - Error
`ifdef SIMULATION
    assert property (@(posedge clk_i) disable iff (!rst_ni)
        mem_if.req_valid |-> can_accept_request)
    else $error("Transaction table overflow detected");

    // AI_TAG: ASSERTION - a_valid_response_opcode: Valid TileLink response opcodes
    assert property (@(posedge clk_i) disable iff (!rst_ni)
        tl_if.d_valid |-> valid_response_opcode)
    else $error("Invalid TileLink response opcode: %h", tl_if.d_opcode);

    // AI_TAG: ASSERTION - a_valid_source_id: Source ID should be within valid range
    assert property (@(posedge clk_i) disable iff (!rst_ni)
        tl_if.a_valid |-> (tl_if.a_source < MAX_OUTSTANDING))
    else $error("Invalid source ID: %d", tl_if.a_source);

    // AI_TAG: ASSERTION - a_valid_response_source_id: Response source ID should match outstanding transaction
    assert property (@(posedge clk_i) disable iff (!rst_ni)
        (tl_if.d_valid && tl_if.d_ready) |-> 
        (transaction_table[tl_if.d_source].valid && 
         transaction_table[tl_if.d_source].tl_source_id == tl_if.d_source))
    else $error("Response source ID does not match outstanding transaction");

    // AI_TAG: ASSERTION - a_tl_req_stable: TileLink request should remain stable when valid
    assert property (@(posedge clk_i) disable iff (!rst_ni)
        tl_if.a_valid && !tl_if.a_ready |=> tl_if.a_valid)
    else $error("TileLink request not stable");
`endif

endmodule : tilelink_adapter

//=============================================================================
// Dependencies: riscv_core_pkg.sv, memory_req_rsp_if.sv, tilelink_if.sv
//
// Performance:
//   - Critical Path: Transaction table lookup and TileLink interface timing
//   - Max Frequency: 500MHz ASIC, 250MHz FPGA
//   - Area: Minimal, optimized for TL-UL subset (~300 gates base + 40 per transaction)
//
// Verification Coverage:
//   - Code Coverage: TBD
//   - Functional Coverage: TileLink protocol compliance
//   - Branch Coverage: All TileLink opcodes and transaction states
//
// Synthesis:
//   - Target Technology: ASIC/FPGA
//   - Synthesis Tool: Design Compiler/Quartus
//   - Clock Domains: 1 (clk_i)
//   - Constraints File: tilelink_adapter.sdc
//
// Testing:
//   - Testbench: tilelink_adapter_tb.sv
//   - Test Vectors: TileLink protocol compliance scenarios
//
//----
// Revision History:
// Version | Date       | Author             | Description
//=============================================================================
// 2.0.0   | 2025-01-27 | DesignAI          | Updated to use proper tilelink_if interface
// 1.0.0   | 2025-01-27 | DesignAI          | Initial TileLink adapter implementation
//============================================================================= 