////////////////////////////////////////////////////////////////////////////////
//
// Company:       Your Company Name
// Engineer:      DesignAI
//
// Create Date:   2025-06-28
// Design Name:   RV32IM Core
// Module Name:   csr_regfile
// Project Name:  riscv_cpu
// Target Devices:ASIC
// Tool Versions:
// Description:   Control and Status Register (CSR) file for the RISC-V core.
//                - Implements essential M-mode CSRs (mstatus, mepc, mcause, etc.).
//                - Handles atomic CSR read/write/set/clear operations from instructions.
//                - Manages state updates during traps (exceptions/interrupts) and mret.
//
// Dependencies:  riscv_core_pkg.sv
//
// Revision:
// Revision 1.0.0 - File Created
// Additional Comments:
//
////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps
`default_nettype none

module csr_regfile
    import riscv_core_pkg::*;
#(
    // AI_TAG: PARAMETER - HART_ID - A unique ID for this processor core (hart).
    parameter word_t HART_ID = 32'd0
)
(
    input  logic        clk_i,
    input  logic        rst_ni,

    // --- CSR Access Port (from Execute stage) ---
    // AI_TAG: PORT_DESC - csr_addr_i - 12-bit address of the CSR to access.
    input  logic [11:0] csr_addr_i,
    // AI_TAG: PORT_DESC - csr_op_i - Type of CSR operation (from funct3: RW, RS, RC).
    input  logic [2:0]  csr_op_i,
    // AI_TAG: PORT_DESC - write_en_i - Asserted for any CSR instruction that writes.
    input  logic        write_en_i,
    // AI_TAG: PORT_DESC - rs1_data_i - Write data operand from rs1 or immediate.
    input  word_t       rs1_data_i,
    // AI_TAG: PORT_DESC - read_data_o - Data read from CSR (value before modification).
    output word_t       read_data_o,

    // --- Trap Control Interface ---
    // AI_TAG: PORT_DESC - trap_en_i - Signals an exception or interrupt is being taken.
    input  logic        trap_en_i,
    // AI_TAG: PORT_DESC - mret_en_i - Signals an MRET instruction is executing.
    input  logic        mret_en_i,
    // AI_TAG: PORT_DESC - mepc_i - PC value to save on a trap.
    input  addr_t       mepc_i,
    // AI_TAG: PORT_DESC - mcause_i - Cause code to save on a trap.
    input  word_t       mcause_i,
    // AI_TAG: PORT_DESC - mtval_i - Trap-specific value (e.g., faulting address).
    input  word_t       mtval_i,

    // --- CSR State Outputs (to control logic) ---
    // AI_TAG: PORT_DESC - mepc_o - Output of MEPC register, used for MRET.
    output addr_t       mepc_o,
    // AI_TAG: PORT_DESC - mtvec_o - Output of MTVEC, the trap vector base address.
    output addr_t       mtvec_o,
    // AI_TAG: PORT_DESC - mstatus_o - Output of MSTATUS register.
    output word_t       mstatus_o
);

    // AI_TAG: RISC-V_SPEC - CSR operation types from instruction's funct3 field.
    localparam logic [2:0] CSR_OP_RW = 3'b001; // CSRRW
    localparam logic [2:0] CSR_OP_RS = 3'b010; // CSRRS
    localparam logic [2:0] CSR_OP_RC = 3'b011; // CSRRC

    // AI_TAG: RISC-V_SPEC - MISA reset value for RV32IM. [31:30]=01 (RV32), [12]=M, [8]=I.
    localparam word_t MISA_RESET_VAL = 32'h40001101;

    // AI_TAG: INTERNAL_STORAGE - Registers for each implemented M-mode CSR.
    word_t mstatus_q, misa_q, mie_q, mtvec_q, mscratch_q, mepc_q, mcause_q, mtval_q, mip_q;
    word_t mhartid_q; // Modeled as a register, but read-only.

    // AI_TAG: INTERNAL_LOGIC - CSR Read Mux
    // Description: Combinational logic to read the current value of a CSR based on its address.
    // This provides the value *before* any modification in the same cycle.
    always_comb begin
        case (csr_addr_i)
            MSTATUS_ADDR:  read_data_o = mstatus_q;
            MISA_ADDR:     read_data_o = misa_q;
            MIE_ADDR:      read_data_o = mie_q;
            MTVEC_ADDR:    read_data_o = mtvec_q;
            MSCRATCH_ADDR: read_data_o = mscratch_q;
            MEPC_ADDR:     read_data_o = mepc_q;
            MCAUSE_ADDR:   read_data_o = mcause_q;
            MTVAL_ADDR:    read_data_o = mtval_q;
            MIP_ADDR:      read_data_o = mip_q;
            MHARTID_ADDR:  read_data_o = mhartid_q;
            default:       read_data_o = '0; // Reads to unimplemented CSRs return 0.
        endcase
    end

    // AI_TAG: INTERNAL_LOGIC - CSR Write and State Update Logic
    // Description: Sequential logic that handles all state changes to the CSRs.
    // Trap handling has the highest priority, followed by MRET, then standard CSR instructions.
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            // Reset values as per RISC-V privileged spec
            mstatus_q  <= '0;
            misa_q     <= MISA_RESET_VAL;
            mie_q      <= '0;
            mtvec_q    <= '0;
            mscratch_q <= '0;
            mepc_q     <= '0;
            mcause_q   <= '0;
            mtval_q    <= '0;
            mip_q      <= '0;
            mhartid_q  <= HART_ID;
        end else begin
            // Priority 1: Trap event (Exception or Interrupt)
            if (trap_en_i) begin
                mepc_q    <= mepc_i;
                mcause_q  <= mcause_i;
                mtval_q   <= mtval_i;
                // Update mstatus: MIE -> MPIE, MIE is cleared
                mstatus_q <= {mstatus_q[31:8], mstatus_q[3], mstatus_q[6:4], 1'b0, mstatus_q[2:0]};
            // Priority 2: MRET instruction
            end else if (mret_en_i) begin
                // Restore previous interrupt-enable state
                mstatus_q <= {mstatus_q[31:8], 1'b1, mstatus_q[6:4], mstatus_q[7], mstatus_q[2:0]};
            // Priority 3: Standard CSR instruction write
            end else if (write_en_i) begin
                case (csr_addr_i)
                    MSTATUS_ADDR:  mstatus_q  <= csr_op(mstatus_q, rs1_data_i, csr_op_i);
                    MIE_ADDR:      mie_q      <= csr_op(mie_q, rs1_data_i, csr_op_i);
                    MTVEC_ADDR:    mtvec_q    <= csr_op(mtvec_q, rs1_data_i, csr_op_i);
                    MSCRATCH_ADDR: mscratch_q <= csr_op(mscratch_q, rs1_data_i, csr_op_i);
                    MEPC_ADDR:     mepc_q     <= csr_op(mepc_q, rs1_data_i, csr_op_i);
                    MCAUSE_ADDR:   mcause_q   <= csr_op(mcause_q, rs1_data_i, csr_op_i);
                    MTVAL_ADDR:    mtval_q    <= csr_op(mtval_q, rs1_data_i, csr_op_i);
                    MIP_ADDR:      mip_q      <= csr_op(mip_q, rs1_data_i, csr_op_i);
                    // MISA and MHARTID are read-only; writes are ignored.
                    default: ;
                endcase
            end
        end
    end

    // AI_TAG: INTERNAL_FUNCTION - csr_op
    // Description: Helper function to perform the atomic CSR operations.
    function automatic word_t csr_op(input word_t csr_val, input word_t write_val, input logic [2:0] op);
        case (op)
            CSR_OP_RW: return write_val;
            CSR_OP_RS: return csr_val | write_val;
            CSR_OP_RC: return csr_val & ~write_val;
            default:   return csr_val; // No operation
        endcase
    endfunction

    // AI_TAG: MODULE_OUTPUTS
    assign mepc_o    = mepc_q;
    assign mtvec_o   = mtvec_q;
    assign mstatus_o = mstatus_q;

endmodule : csr_regfile

`default_nettype wire