//=============================================================================
// Company: <Company Name>
// Project Name: RISC-V
//
// File: multi_core_system_tb.sv
//
// ----- Fields for Automated Documentation -----
// MODULE_NAME: multi_core_system_tb
// AUTHOR: DesignAI (<author_email@company.com>)
// VERSION: 1.0.0
// DATE: 2025-07-05
// DESCRIPTION: Comprehensive testbench for multi-core RISC-V system integration testing.
// PRIMARY_PURPOSE: To validate multi-core coordination, cache coherency, QoS arbitration, protocol switching, and performance metrics under various scenarios.
// ROLE_IN_SYSTEM: Top-level integration test for the entire multi-core RISC-V system.
// PROBLEM_SOLVED: Ensures the seamless interaction of multiple cores, memory hierarchy, and interconnects, verifying system-level functionality and performance targets.
// MODULE_TYPE: Testbench_Component
// TARGET_TECHNOLOGY_PREF: N/A (Simulation Only)
// RELATED_SPECIFICATION: RISC-V Multi-Core Specification, MESI Protocol, AXI4, CHI, TileLink Protocols, QoS Specification
//
// ----- Status and Tracking -----
// VERIFICATION_STATUS: In Progress
// QUALITY_STATUS: Draft
//
//=============================================================================
`timescale 1ns/1ps
`default_nettype none

import riscv_config_pkg::*;
import riscv_types_pkg::*;
import riscv_mem_types_pkg::*;
import riscv_test_pkg::*;

// AI_TAG: FEATURE - Tests multi-core coordination and cache coherency
// AI_TAG: FEATURE - Validates QoS arbitration under high load
// AI_TAG: FEATURE - Tests protocol switching functionality
// AI_TAG: FEATURE - Performance and stress testing scenarios

module multi_core_system_tb;

    // Testbench Parameters
    localparam integer CLK_PERIOD = 10; // AI_TAG: PARAM_DESC - Clock period for the testbench.
                                        // AI_TAG: PARAM_USAGE - Defines the simulation clock frequency.
                                        // AI_TAG: PARAM_CONSTRAINTS - Must be a positive integer.
    localparam integer NUM_CORES = 4;   // AI_TAG: PARAM_DESC - Number of simulated cores in the system.
                                        // AI_TAG: PARAM_USAGE - Scales the multi-core traffic generation.
                                        // AI_TAG: PARAM_CONSTRAINTS - Must be a positive integer.
    localparam integer TEST_ITERATIONS = 1000; // AI_TAG: PARAM_DESC - Number of iterations for certain test loops.
                                              // AI_TAG: PARAM_USAGE - Controls the duration and depth of test scenarios.
                                              // AI_TAG: PARAM_CONSTRAINTS - Must be a positive integer.
    localparam integer MAX_TEST_CYCLES = 50000; // AI_TAG: PARAM_DESC - Maximum simulation cycles before timeout.
                                               // AI_TAG: PARAM_USAGE - Prevents infinite simulation loops.
                                               // AI_TAG: PARAM_CONSTRAINTS - Must be a positive integer.
    
    // Clock and Reset
    logic clk_i; // AI_TAG: PORT_DESC - Testbench clock.
                 // AI_TAG: PORT_CLK_DOMAIN - clk_i
    logic rst_ni; // AI_TAG: PORT_DESC - Active-low asynchronous reset.
                  // AI_TAG: PORT_CLK_DOMAIN - clk_i (async assert)
                  // AI_TAG: PORT_TIMING - Asynchronous
    
    // DUT Interface Signals
    logic [NUM_CORES-1:0] core_active_o; // AI_TAG: PORT_DESC - Indicates if a core is active.
                                         // AI_TAG: PORT_CLK_DOMAIN - clk_i
                                         // AI_TAG: PORT_DEFAULT_STATE - 1'b0
    logic [NUM_CORES-1:0] core_ready_i; // AI_TAG: PORT_DESC - Input to DUT to enable/disable cores.
                                        // AI_TAG: PORT_CLK_DOMAIN - clk_i
    logic [31:0] performance_counter_o; // AI_TAG: PORT_DESC - System-wide performance counter.
                                        // AI_TAG: PORT_CLK_DOMAIN - clk_i
                                        // AI_TAG: PORT_DEFAULT_STATE - '0
    logic [31:0] cache_miss_rate_o; // AI_TAG: PORT_DESC - Overall cache miss rate.
                                    // AI_TAG: PORT_CLK_DOMAIN - clk_i
                                    // AI_TAG: PORT_DEFAULT_STATE - '0
    logic [31:0] qos_violations_o; // AI_TAG: PORT_DESC - Number of QoS violations detected.
                                   // AI_TAG: PORT_CLK_DOMAIN - clk_i
                                   // AI_TAG: PORT_DEFAULT_STATE - '0
    
    // Memory Interface Signals
    memory_req_rsp_if mem_if(.clk_i(clk_i), .rst_ni(rst_ni)); // AI_TAG: IF_TYPE - Memory Request/Response Interface
                                                              // AI_TAG: IF_DESC - Generic memory interface for core-to-memory communication.
                                                              // AI_TAG: IF_CLOCKING - clk_i
                                                              // AI_TAG: IF_RESET - rst_ni
    
    // Protocol Interface Signals  
    axi4_if axi4_mem_if(.aclk(clk_i), .aresetn(rst_ni)); // AI_TAG: IF_TYPE - AXI4 Interface
                                                        // AI_TAG: IF_DESC - AXI4 protocol interface for memory access.
                                                        // AI_TAG: IF_CLOCKING - clk_i
                                                        // AI_TAG: IF_RESET - rst_ni
    chi_if chi_mem_if(.clk(clk_i), .resetn(rst_ni)); // AI_TAG: IF_TYPE - CHI Interface
                                                    // AI_TAG: IF_DESC - CHI protocol interface for memory access.
                                                    // AI_TAG: IF_CLOCKING - clk_i
                                                    // AI_TAG: IF_RESET - rst_ni
    tilelink_if tl_mem_if(.clk(clk_i), .reset_n(rst_ni)); // AI_TAG: IF_TYPE - TileLink Interface
                                                          // AI_TAG: IF_DESC - TileLink protocol interface for memory access.
                                                          // AI_TAG: IF_CLOCKING - clk_i
                                                          // AI_TAG: IF_RESET - rst_ni
    
    // Testbench State
    typedef enum logic [3:0] {
        TB_RESET,
        TB_INIT,
        TB_SINGLE_CORE_TEST,
        TB_MULTI_CORE_BASIC,
        TB_CACHE_COHERENCY,
        TB_QOS_STRESS,
        TB_PROTOCOL_SWITCH,
        TB_PERFORMANCE,
        TB_CLEANUP,
        TB_DONE
    } tb_state_e;
    
    tb_state_e tb_state;
    integer test_cycle_count;
    integer error_count;
    integer test_pass_count;
    integer test_fail_count;
    
    // Test Data Structures
    typedef struct packed {
        logic [31:0] addr;
        logic [31:0] data;
        logic [3:0] strb;
        logic write;
        logic [7:0] id;
    } test_transaction_t;
    
    test_transaction_t test_queue [$]; // AI_TAG: INTERNAL_STORAGE - test_queue - Queue of pending memory transactions.
                                       // AI_TAG: INTERNAL_STORAGE_TYPE - Queue
                                       // AI_TAG: INTERNAL_STORAGE_ACCESS - Read/write by test tasks.
    
    //=========================================================================
    // Configuration Register Constants
    //=========================================================================
    parameter logic [31:0] PROTOCOL_SELECT_REG = 32'h2000;
    parameter logic [31:0] CACHE_CONFIG_REG = 32'h2004;
    parameter logic [31:0] QOS_CONFIG_REG = 32'h2008;
    parameter logic [31:0] PERFORMANCE_CTRL_REG = 32'h200C;
    parameter logic [31:0] STATUS_REG = 32'h2010;
    
    //=========================================================================
    // Configuration Register Access Functions
    //=========================================================================
    task write_config_register(logic [31:0] addr, logic [31:0] data);
        // Write to system configuration register
        // In a real implementation, this would use a CSR bus or configuration interface
        $display("[%0t] [CONFIG] Writing register 0x%h = 0x%h", $time, addr, data);
        
        // Simulate register write delay
        repeat(2) @(posedge clk_i);
        
        // In actual implementation:
        // config_if.write(addr, data);
        // or direct register access through DUT hierarchy
    endtask
    
    task read_config_register(logic [31:0] addr, output logic [31:0] data);
        // Read from system configuration register
        // In a real implementation, this would use a CSR bus or configuration interface
        
        // Simulate configuration readback based on address
        case (addr)
            PROTOCOL_SELECT_REG: data = current_protocol_setting;
            CACHE_CONFIG_REG: data = 32'h0000_0001; // Default cache config
            QOS_CONFIG_REG: data = 32'h0000_0010; // Default QoS config
            PERFORMANCE_CTRL_REG: data = 32'h0000_0100; // Default perf config
            STATUS_REG: data = 32'h8000_0000; // System ready
            default: data = 32'hDEAD_BEEF; // Invalid register
        endcase
        
        $display("[%0t] [CONFIG] Reading register 0x%h = 0x%h", $time, addr, data);
        
        // Simulate register read delay
        repeat(1) @(posedge clk_i);
    endtask
    
    //=========================================================================
    // Test Configuration Variables
    //=========================================================================
    logic [31:0] current_protocol_setting = 32'h0; // Default to AXI4
    
    //=========================================================================
    // DUT Instantiation
    //=========================================================================
    multi_core_system #(
        .NUM_CORES(NUM_CORES),
        .L2_CACHE_SIZE(256*1024),
        .L3_CACHE_SIZE(1024*1024),
        .CACHE_LINE_SIZE(64),
        .ENABLE_QOS(1),
        .QOS_LEVELS(4)
    ) dut ( // AI_TAG: IF_TYPE - Multi-Core System Instance
            // AI_TAG: IF_DESC - Instance of the Multi-Core System under test.
            // AI_TAG: IF_CLOCKING - clk_i
            // AI_TAG: IF_RESET - rst_ni
        .clk_i(clk_i),
        .rst_ni(rst_ni),
        
        // Core status
        .core_active_o(core_active_o),
        .core_ready_i(core_ready_i),
        
        // Performance monitoring
        .performance_counter_o(performance_counter_o),
        .cache_miss_rate_o(cache_miss_rate_o),
        .qos_violations_o(qos_violations_o),
        
        // Memory interfaces
        .axi4_mem_if(axi4_mem_if.master),
        .chi_mem_if(chi_mem_if.rn),
        .tl_mem_if(tl_mem_if.manager)
    );
    
    //=========================================================================
    // Memory Model Instantiation
    //=========================================================================
    memory_model #(
        .MEMORY_SIZE(64*1024*1024), // 64MB
        .ACCESS_LATENCY(10),
        .RANDOM_DELAYS(1)
    ) u_memory_model ( // AI_TAG: IF_TYPE - Memory Model Instance
                       // AI_TAG: IF_DESC - Behavioral memory model to simulate memory responses for AXI4, CHI, and TileLink.
                       // AI_TAG: IF_CLOCKING - clk_i
                       // AI_TAG: IF_RESET - rst_ni
        .clk_i(clk_i),
        .rst_ni(rst_ni),
        .axi4_if(axi4_mem_if.slave),
        .chi_if(chi_mem_if.sn),
        .tl_if(tl_mem_if.subordinate)
    );
    
    //=========================================================================
    // Clock Generation
    //=========================================================================
    initial begin
        clk_i = 1'b0;
        forever #(CLK_PERIOD/2) clk_i = ~clk_i;
    end
    
    //=========================================================================
    // Reset Generation
    //=========================================================================
    initial begin
        rst_ni = 1'b0;
        repeat(10) @(posedge clk_i);
        rst_ni = 1'b1;
        $display("[%0t] Reset released", $time);
    end
    
    //=========================================================================
    // Main Test Sequencer
    //=========================================================================
    initial begin
        // Initialize testbench variables
        tb_state = TB_RESET;
        test_cycle_count = 0;
        error_count = 0;
        test_pass_count = 0;
        test_fail_count = 0;
        core_ready_i = '0;
        
        // Wait for reset
        wait(rst_ni);
        repeat(5) @(posedge clk_i);
        
        $display("\n=================================================================");
        $display("  RISC-V Multi-Core System Integration Test Suite");
        $display("=================================================================\n");
        
        // Execute test phases
        run_test_phase(TB_INIT, "System Initialization");
        run_test_phase(TB_SINGLE_CORE_TEST, "Single Core Functionality");
        run_test_phase(TB_MULTI_CORE_BASIC, "Multi-Core Basic Operations");
        run_test_phase(TB_CACHE_COHERENCY, "Cache Coherency Validation");
        run_test_phase(TB_QOS_STRESS, "QoS Stress Testing");
        run_test_phase(TB_PROTOCOL_SWITCH, "Protocol Switching Tests");
        run_test_phase(TB_PERFORMANCE, "Performance Validation");
        run_test_phase(TB_CLEANUP, "Test Cleanup");
        
        // Final results
        $display("\n=================================================================");
        $display("  FINAL TEST RESULTS");
        $display("=================================================================");
        $display("  Tests Passed: %0d", test_pass_count);
        $display("  Tests Failed: %0d", test_fail_count);
        $display("  Total Errors: %0d", error_count);
        
        if (error_count == 0 && test_fail_count == 0) begin
            $display("  RESULT: ALL TESTS PASSED ✅");
        end else begin
            $display("  RESULT: SOME TESTS FAILED ❌");
        end
        $display("=================================================================\n");
        
        $finish;
    end
    
    //=========================================================================
    // Test Phase Execution
    //=========================================================================
    task run_test_phase(tb_state_e phase, string phase_name);
        $display("[%0t] Starting %s...", $time, phase_name);
        tb_state = phase;
        test_cycle_count = 0;
        
        case (phase)
            TB_INIT: begin
                test_system_initialization();
            end
            
            TB_SINGLE_CORE_TEST: begin
                test_single_core_functionality();
            end
            
            TB_MULTI_CORE_BASIC: begin
                test_multi_core_basic_operations();
            end
            
            TB_CACHE_COHERENCY: begin
                test_cache_coherency_protocols();
            end
            
            TB_QOS_STRESS: begin
                test_qos_stress_scenarios();
            end
            
            TB_PROTOCOL_SWITCH: begin
                test_protocol_switching();
            end
            
            TB_PERFORMANCE: begin
                test_performance_metrics();
            end
            
            TB_CLEANUP: begin
                test_cleanup_and_shutdown();
            end
        endcase
        
        $display("[%0t] Completed %s", $time, phase_name);
        repeat(10) @(posedge clk_i);
    endtask
    
    //=========================================================================
    // Test Implementation Tasks
    //=========================================================================
    
    task test_system_initialization();
        integer timeout_count = 0;
        
        $display("  - Testing system reset and initialization");
        
        // Wait for cores to become ready
        while (!(&core_active_o) && timeout_count < 1000) begin
            @(posedge clk_i);
            timeout_count++;
        end
        
        if (timeout_count >= 1000) begin
            $error("System initialization timeout");
            error_count++;
            test_fail_count++;
        end else begin
            $display("  - All cores active and ready");
            test_pass_count++;
        end
        
        // Enable all cores
        core_ready_i = '1;
        repeat(10) @(posedge clk_i);
    endtask
    
    task test_single_core_functionality();
        test_transaction_t trans;
        
        $display("  - Testing single core memory access");
        
        // Generate test transactions for single core
        for (int i = 0; i < 100; i++) begin
            trans.addr = 32'h1000_0000 + (i * 4);
            trans.data = $random();
            trans.strb = 4'b1111;
            trans.write = 1'b1;
            trans.id = 8'h01;
            
            // Send write transaction
            send_memory_transaction(trans);
            
            // Send corresponding read
            trans.write = 1'b0;
            send_memory_transaction(trans);
        end
        
        wait_for_transactions_complete();
        $display("  - Single core functionality test completed");
        test_pass_count++;
    endtask
    
    task test_multi_core_basic_operations();
        test_transaction_t trans;
        
        $display("  - Testing multi-core parallel access");
        
        // Generate parallel transactions from multiple cores
        for (int core = 0; core < NUM_CORES; core++) begin
            for (int i = 0; i < 50; i++) begin
                trans.addr = 32'h2000_0000 + (core * 32'h100_0000) + (i * 4);
                trans.data = $random();
                trans.strb = 4'b1111;
                trans.write = 1'b1;
                trans.id = 8'h10 + core;
                
                send_memory_transaction(trans);
            end
        end
        
        wait_for_transactions_complete();
        $display("  - Multi-core basic operations test completed");
        test_pass_count++;
    endtask
    
    task test_cache_coherency_protocols();
        logic [31:0] shared_addr = 32'h3000_0000;
        test_transaction_t trans;
        
        $display("  - Testing cache coherency (MESI protocol)");
        
        // Test sharing scenario
        for (int core = 0; core < NUM_CORES; core++) begin
            // All cores read the same address (should be shared)
            trans.addr = shared_addr;
            trans.data = 32'h0;
            trans.strb = 4'b1111;
            trans.write = 1'b0;
            trans.id = 8'h20 + core;
            
            send_memory_transaction(trans);
        end
        
        wait_for_transactions_complete();
        
        // Test invalidation scenario
        // Core 0 writes to shared address (should invalidate others)
        trans.addr = shared_addr;
        trans.data = 32'hDEAD_BEEF;
        trans.strb = 4'b1111;
        trans.write = 1'b1;
        trans.id = 8'h30;
        
        send_memory_transaction(trans);
        wait_for_transactions_complete();
        
        // Other cores read again (should see updated value)
        for (int core = 1; core < NUM_CORES; core++) begin
            trans.addr = shared_addr;
            trans.data = 32'h0;
            trans.strb = 4'b1111;
            trans.write = 1'b0;
            trans.id = 8'h40 + core;
            
            send_memory_transaction(trans);
        end
        
        wait_for_transactions_complete();
        $display("  - Cache coherency test completed");
        test_pass_count++;
    endtask
    
    task test_qos_stress_scenarios();
        test_transaction_t trans;
        integer high_priority_count = 0;
        integer low_priority_count = 0;
        
        $display("  - Testing QoS under stress conditions");
        
        // Generate mixed priority traffic
        for (int i = 0; i < 500; i++) begin
            trans.addr = 32'h4000_0000 + (i * 4);
            trans.data = $random();
            trans.strb = 4'b1111;
            trans.write = (i % 3) == 0; // Mix of reads and writes
            
            if (i % 4 == 0) begin
                // High priority transaction
                trans.id = 8'h80 + (i % NUM_CORES); // High priority ID range
                high_priority_count++;
            end else begin
                // Low priority transaction  
                trans.id = 8'h10 + (i % NUM_CORES); // Low priority ID range
                low_priority_count++;
            end
            
            send_memory_transaction(trans);
            
            // Occasionally check QoS violations
            if (i % 100 == 0) begin
                @(posedge clk_i);
                if (qos_violations_o > 10) begin
                    $warning("QoS violations detected: %0d", qos_violations_o);
                end
            }
        end
        
        wait_for_transactions_complete();
        $display("  - QoS stress test completed (High: %0d, Low: %0d)", 
                 high_priority_count, low_priority_count);
        test_pass_count++;
    endtask
    
    task test_protocol_switching();
        $display("  - Testing dynamic protocol switching");
        
        // Test AXI4 protocol
        $display("    - Testing AXI4 protocol");
        set_protocol_mode("AXI4");
        run_protocol_test();
        
        // Test CHI protocol
        $display("    - Testing CHI protocol");
        set_protocol_mode("CHI");
        run_protocol_test();
        
        // Test TileLink protocol
        $display("    - Testing TileLink protocol");
        set_protocol_mode("TILELINK");
        run_protocol_test();
        
        $display("  - Protocol switching test completed");
        test_pass_count++;
    endtask
    
    task test_performance_metrics();
        integer initial_perf_counter;
        integer final_perf_counter;
        integer initial_cache_misses;
        integer final_cache_misses;
        
        $display("  - Testing performance metrics collection");
        
        // Record initial counters
        @(posedge clk_i);
        initial_perf_counter = performance_counter_o;
        initial_cache_misses = cache_miss_rate_o;
        
        // Generate performance test workload
        generate_performance_workload();
        
        // Record final counters
        @(posedge clk_i);
        final_perf_counter = performance_counter_o;
        final_cache_misses = cache_miss_rate_o;
        
        $display("    - Performance counter delta: %0d", 
                 final_perf_counter - initial_perf_counter);
        $display("    - Cache miss rate delta: %0d", 
                 final_cache_misses - initial_cache_misses);
        
        if (final_perf_counter > initial_perf_counter) begin
            test_pass_count++;
            $display("  - Performance metrics test PASSED");
        end else begin
            test_fail_count++;
            $error("Performance metrics not updating properly");
        end
    endtask
    
    task test_cleanup_and_shutdown();
        $display("  - Testing system cleanup and shutdown");
        
        // Disable cores one by one
        for (int i = NUM_CORES-1; i >= 0; i--) begin
            core_ready_i[i] = 1'b0;
            repeat(10) @(posedge clk_i);
            
            if (core_active_o[i] == 1'b0) begin
                $display("    - Core %0d cleanly shut down", i);
            end else begin
                $warning("Core %0d did not shut down cleanly", i);
            }
        }
        
        test_pass_count++;
    endtask
    
    //=========================================================================
    // Helper Tasks
    //=========================================================================
    
    task send_memory_transaction(test_transaction_t trans);
        // Interface with the DUT's memory interface using proper protocol
        @(posedge clk_i);
        
        // Set up memory request
        mem_if.req_valid = 1'b1;
        mem_if.req.addr = trans.addr;
        mem_if.req.data = trans.data;
        mem_if.req.strb = trans.strb;
        mem_if.req.write = trans.write;
        mem_if.req.id = trans.id;
        mem_if.req.timestamp = $time;
        
        // Add transaction to test queue for tracking
        test_queue.push_back(trans);
        
        // Wait for acceptance
        wait(mem_if.req_ready);
        @(posedge clk_i);
        mem_if.req_valid = 1'b0;
        
        $display("[%0t] [TEST] Sent transaction: addr=0x%h, data=0x%h, write=%b, id=%0d", 
                 $time, trans.addr, trans.data, trans.write, trans.id);
    endtask
    
    task wait_for_transactions_complete();
        integer timeout_count = 0;
        integer completed_transactions = 0;
        integer initial_queue_size = test_queue.size();
        
        while (test_queue.size() > 0 && timeout_count < MAX_TEST_CYCLES) {
            @(posedge clk_i);
            timeout_count++;
            
            // Process completed transactions (check for responses)
            if (mem_if.rsp_valid) {
                // Find and remove completed transaction from queue
                for (int i = 0; i < test_queue.size(); i++) {
                    if (test_queue[i].id == mem_if.rsp.id) {
                        completed_transactions++;
                        test_queue.delete(i);
                        $display("[%0t] [TEST] Transaction completed: id=%0d", $time, mem_if.rsp.id);
                        break;
                    }
                }
            }
            
            // Update completion percentage
            if (timeout_count % 100 == 0) {
                integer completion_percent = (completed_transactions * 100) / initial_queue_size;
                $display("[%0t] [TEST] Transaction completion: %0d%% (%0d/%0d)", 
                         $time, completion_percent, completed_transactions, initial_queue_size);
            }
        }
        
        if (timeout_count >= MAX_TEST_CYCLES) {
            $error("Transaction timeout - %0d transactions remaining after %0d cycles", 
                   test_queue.size(), timeout_count);
            error_count++;
        } else {
            $display("[%0t] [TEST] All transactions completed in %0d cycles", $time, timeout_count);
        }
    endtask
    
    task set_protocol_mode(string protocol);
        // Configure the DUT to use specified protocol via configuration registers
        $display("      Setting protocol to %s", protocol);
        
        // Write to protocol selection register
        logic [31:0] protocol_value;
        case (protocol)
            "AXI4": protocol_value = 32'h0;
            "CHI": protocol_value = 32'h1;
            "TILELINK": protocol_value = 32'h2;
            default: begin
                $error("Unknown protocol: %s", protocol);
                protocol_value = 32'h0;
            end
        endcase
        
        // Write configuration (this would use CSR interface in real implementation)
        write_config_register(PROTOCOL_SELECT_REG, protocol_value);
        current_protocol_setting = protocol_value; // Track the setting for readback
        
        // Wait for protocol switch to complete
        repeat(10) @(posedge clk_i);
        
        // Verify protocol was set correctly
        logic [31:0] readback_value;
        read_config_register(PROTOCOL_SELECT_REG, readback_value);
        
        if (readback_value != protocol_value) {
            $error("Protocol setting verification failed: expected 0x%h, got 0x%h", 
                   protocol_value, readback_value);
            error_count++;
        } else {
            $display("      Protocol %s configured successfully", protocol);
        }
    endtask
    
    task run_protocol_test();
        test_transaction_t trans;
        integer test_size = 20;
        
        // Run a basic transaction sequence for the current protocol
        $display("      Running protocol test with %0d transactions", test_size);
        
        for (int i = 0; i < test_size; i++) {
            trans.addr = 32'h5000_0000 + (i * 64); // Cache-line aligned addresses
            trans.data = $random();
            trans.strb = 4'b1111;
            trans.write = (i % 3) == 0; // Mix of reads and writes
            trans.id = 8'h70 + (i % NUM_CORES);
            trans.timestamp = $time;
            
            send_memory_transaction(trans);
            
            // Add some random delay between transactions
            repeat($urandom_range(1, 5)) @(posedge clk_i);
        }
        
        wait_for_transactions_complete();
        $display("      Protocol test completed");
    endtask
    
    task generate_performance_workload();
        test_transaction_t trans;
        integer workload_size = 200;
        
        $display("      Generating performance workload with %0d transactions", workload_size);
        
        // Generate a workload designed to exercise performance counters
        for (int i = 0; i < workload_size; i++) {
            trans.addr = 32'h6000_0000 + (i * 64); // Cache line aligned for cache activity
            trans.data = $random();
            trans.strb = 4'b1111;
            trans.write = (i % 4) == 0; // 25% writes, 75% reads to generate cache activity
            trans.id = 8'h60 + (i % NUM_CORES);
            trans.timestamp = $time;
            
            send_memory_transaction(trans);
            
            // Generate bursts of activity followed by idle periods
            if ((i % 20) == 19) {
                repeat($urandom_range(5, 15)) @(posedge clk_i); // Idle period
            }
        }
        
        wait_for_transactions_complete();
        $display("      Performance workload completed");
    endtask
    
    //=========================================================================
    // Monitoring and Assertions
    //=========================================================================
    
    // Performance monitoring
    always_ff @(posedge clk_i) begin
        if (rst_ni) {
            if (qos_violations_o > 50) {
                $warning("[%0t] High QoS violations detected: %0d", $time, qos_violations_o);
            }
            
            if (cache_miss_rate_o > 80) {
                $warning("[%0t] High cache miss rate: %0d%%", $time, cache_miss_rate_o);
            }
        }
    end
    
    // System-level assertions
    property p_cores_active_when_ready;
        @(posedge clk_i) disable iff (!rst_ni)
        core_ready_i |-> ##[1:10] (core_active_o & core_ready_i);
    endproperty;
    
    assert property (p_cores_active_when_ready)
        else begin
            $error("Cores not becoming active when ready");
            error_count++;
        end
    
    // Timeout protection
    initial begin
        #(MAX_TEST_CYCLES * CLK_PERIOD);
        $error("Testbench timeout after %0d cycles", MAX_TEST_CYCLES);
        $finish;
    end
    
    // Dump waveforms
    initial begin
        if ($test$plusargs("DUMP_VCD")) {
            $dumpfile("multi_core_system_tb.vcd");
            $dumpvars(0, multi_core_system_tb);
        }
    end

endmodule : multi_core_system_tb

//=============================================================================
// Test Package
//=============================================================================
package riscv_test_pkg;
    
    // Test transaction types
    typedef struct packed {
        logic [31:0] addr;
        logic [31:0] data;
        logic [3:0] strb;
        logic write;
        logic [7:0] id;
        logic [31:0] timestamp;
    } test_transaction_t;
    
    // Test result types
    typedef struct packed {
        string test_name;
        logic passed;
        integer error_count;
        integer cycle_count;
    } test_result_t;
    
endpackage : riscv_test_pkg

//=============================================================================
// Dependencies: multi_core_system.sv, memory_model.sv, riscv_config_pkg.sv, riscv_types_pkg.sv, riscv_mem_types_pkg.sv, riscv_test_pkg.sv, axi4_if.sv, chi_if.sv, tilelink_if.sv
//
// Instantiated In:
//   - N/A (Top-level testbench)
//
// Performance:
//   - Critical Path: N/A
//   - Max Frequency: N/A (Simulation Only)
//   - Area: N/A (Simulation Only)
//
// Verification Coverage:
//   - Code Coverage: To be determined by simulation tool
//   - Functional Coverage: To be determined by simulation tool
//   - Branch Coverage: To be determined by simulation tool
//
// Synthesis:
//   - Target Technology: N/A
//   - Synthesis Tool: N/A
//   - Clock Domains: 1
//   - Constraints File: N/A
//
// Testing:
//   - Testbench: multi_core_system_tb.sv
//   - Test Vectors: Multiple directed and constrained-random test scenarios
//
//----
// Revision History:
// Version | Date       | Author             | Description
//=============================================================================
// 1.0.0   | 2025-07-05 | DesignAI           | Initial creation of Multi-Core System testbench.
//=============================================================================