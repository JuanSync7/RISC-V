////////////////////////////////////////////////////////////////////////////////
//
// Testbench:    icache_tb
// Description:  Unit testbench for the ICache module
//
////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps
`default_nettype none

module icache_tb;
    import riscv_core_pkg::*;

    // Parameters
    localparam CACHE_SIZE = 4096;
    localparam LINE_SIZE  = 32;
    localparam WAYS       = 2;
    localparam ADDR_WIDTH = 32;
    localparam XLEN       = 32;

    // Clock and reset
    logic clk;
    logic rst_n;

    // ICache interface signals
    logic        valid_i;
    addr_t       pc_i;
    logic        ready_o;
    word_t       instruction_o;
    logic        hit_o;
    logic        valid_o;
    // Memory interface
    logic        mem_arvalid_o;
    logic        mem_arready_i;
    addr_t       mem_araddr_o;
    logic        mem_rvalid_i;
    word_t       mem_rdata_i;
    logic        mem_rready_o;
    // Control
    logic        flush_i;
    logic        flush_done_o;

    // Instantiate ICache
    icache #(
        .CACHE_SIZE(CACHE_SIZE),
        .LINE_SIZE(LINE_SIZE),
        .WAYS(WAYS)
    ) dut (
        .clk_i(clk),
        .rst_ni(rst_n),
        .pc_i(pc_i),
        .valid_i(valid_i),
        .ready_o(ready_o),
        .instruction_o(instruction_o),
        .hit_o(hit_o),
        .valid_o(valid_o),
        .mem_arvalid_o(mem_arvalid_o),
        .mem_arready_i(mem_arready_i),
        .mem_araddr_o(mem_araddr_o),
        .mem_rvalid_i(mem_rvalid_i),
        .mem_rdata_i(mem_rdata_i),
        .mem_rready_o(mem_rready_o),
        .flush_i(flush_i),
        .flush_done_o(flush_done_o)
    );

    // Clock generation
    initial clk = 0;
    always #5 clk = ~clk;

    // Test stimulus
    initial begin
        rst_n = 0;
        valid_i = 0;
        pc_i = 0;
        mem_arready_i = 0;
        mem_rvalid_i = 0;
        mem_rdata_i = 0;
        flush_i = 0;
        #20;
        rst_n = 1;
        #10;

        // Test 1: Simple miss and fill
        $display("[TB] Test 1: Simple miss and fill");
        pc_i = 32'h0000_0000;
        valid_i = 1;
        @(posedge clk);
        valid_i = 0;
        // Wait for cache miss and memory request
        wait (mem_arvalid_o);
        $display("[TB] Cache miss detected, memory request issued at addr %h", mem_araddr_o);
        mem_arready_i = 1;
        @(posedge clk);
        mem_arready_i = 0;
        // Simulate memory returning data for the whole line
        repeat (LINE_SIZE/4) begin
            mem_rvalid_i = 1;
            mem_rdata_i = $random;
            @(posedge clk);
        end
        mem_rvalid_i = 0;
        // Wait for cache to become ready
        wait (ready_o);
        $display("[TB] Cache line filled, ready for next request");
        // Issue the same request again (should be a hit)
        valid_i = 1;
        @(posedge clk);
        valid_i = 0;
        @(posedge clk);
        if (hit_o && valid_o)
            $display("[TB] Cache hit for addr %h, instruction: %h", pc_i, instruction_o);
        else
            $display("[TB] ERROR: Expected cache hit");

        // Test 2: Cache flush
        $display("[TB] Test 2: Cache flush");
        flush_i = 1;
        @(posedge clk);
        flush_i = 0;
        wait (flush_done_o);
        $display("[TB] Cache flush done");
        // Issue the same request again (should be a miss)
        valid_i = 1;
        @(posedge clk);
        valid_i = 0;
        wait (mem_arvalid_o);
        $display("[TB] Cache miss after flush as expected");
        mem_arready_i = 1;
        repeat (LINE_SIZE/4) begin
            mem_rvalid_i = 1;
            mem_rdata_i = $random;
            @(posedge clk);
        end
        mem_rvalid_i = 0;
        mem_arready_i = 0;
        wait (ready_o);
        $display("[TB] Cache line refilled after flush");

        // Test 3: LRU Replacement Policy
        $display("[TB] Test 3: LRU Replacement Policy");
        // Access two addresses mapping to the same set but different ways
        logic [31:0] set_base = 32'h1000_0000;
        logic [31:0] addr_a = set_base;
        logic [31:0] addr_b = set_base | (1 << (ADDR_WIDTH-1)); // Different tag, same set
        logic [31:0] addr_c = set_base | (2 << (ADDR_WIDTH-1)); // Third tag, same set
        // Fill way 0
        pc_i = addr_a;
        valid_i = 1;
        @(posedge clk); valid_i = 0;
        wait (mem_arvalid_o); mem_arready_i = 1; @(posedge clk); mem_arready_i = 0;
        repeat (LINE_SIZE/4) begin mem_rvalid_i = 1; mem_rdata_i = $random; @(posedge clk); end
        mem_rvalid_i = 0; wait (ready_o);
        // Fill way 1
        pc_i = addr_b;
        valid_i = 1;
        @(posedge clk); valid_i = 0;
        wait (mem_arvalid_o); mem_arready_i = 1; @(posedge clk); mem_arready_i = 0;
        repeat (LINE_SIZE/4) begin mem_rvalid_i = 1; mem_rdata_i = $random; @(posedge clk); end
        mem_rvalid_i = 0; wait (ready_o);
        // Both should be hits
        pc_i = addr_a; valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
        if (hit_o && valid_o) $display("[TB] LRU: Hit way 0 as expected"); else $display("[TB] ERROR: LRU: Miss on way 0");
        pc_i = addr_b; valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
        if (hit_o && valid_o) $display("[TB] LRU: Hit way 1 as expected"); else $display("[TB] ERROR: LRU: Miss on way 1");
        // Access a third address mapping to same set (should evict LRU)
        pc_i = addr_c; valid_i = 1; @(posedge clk); valid_i = 0;
        wait (mem_arvalid_o); mem_arready_i = 1; @(posedge clk); mem_arready_i = 0;
        repeat (LINE_SIZE/4) begin mem_rvalid_i = 1; mem_rdata_i = $random; @(posedge clk); end
        mem_rvalid_i = 0; wait (ready_o);
        // Now, one of addr_a or addr_b should be evicted (LRU)
        pc_i = addr_a; valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
        if (hit_o && valid_o) $display("[TB] LRU: addr_a still present (expected if addr_b was LRU)");
        else $display("[TB] LRU: addr_a evicted (expected if it was LRU)");
        pc_i = addr_b; valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
        if (hit_o && valid_o) $display("[TB] LRU: addr_b still present (expected if addr_a was LRU)");
        else $display("[TB] LRU: addr_b evicted (expected if it was LRU)");
        pc_i = addr_c; valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
        if (hit_o && valid_o) $display("[TB] LRU: addr_c present as expected");
        else $display("[TB] ERROR: LRU: addr_c not present");

        // Test 4: Associativity (two addresses in same set, both present)
        $display("[TB] Test 4: Associativity");
        // Already covered in Test 3, but repeat for clarity
        pc_i = addr_a; valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
        if (hit_o && valid_o) $display("[TB] Associativity: addr_a hit");
        else $display("[TB] ERROR: Associativity: addr_a miss");
        pc_i = addr_b; valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
        if (hit_o && valid_o) $display("[TB] Associativity: addr_b hit");
        else $display("[TB] ERROR: Associativity: addr_b miss");

        // Test 5: Multiple sets (addresses in different sets, no interference)
        $display("[TB] Test 5: Multiple sets");
        logic [31:0] set2_base = 32'h2000_0000;
        logic [31:0] set3_base = 32'h3000_0000;
        pc_i = set2_base; valid_i = 1; @(posedge clk); valid_i = 0;
        wait (mem_arvalid_o); mem_arready_i = 1; @(posedge clk); mem_arready_i = 0;
        repeat (LINE_SIZE/4) begin mem_rvalid_i = 1; mem_rdata_i = $random; @(posedge clk); end
        mem_rvalid_i = 0; wait (ready_o);
        pc_i = set3_base; valid_i = 1; @(posedge clk); valid_i = 0;
        wait (mem_arvalid_o); mem_arready_i = 1; @(posedge clk); mem_arready_i = 0;
        repeat (LINE_SIZE/4) begin mem_rvalid_i = 1; mem_rdata_i = $random; @(posedge clk); end
        mem_rvalid_i = 0; wait (ready_o);
        // Both should be hits
        pc_i = set2_base; valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
        if (hit_o && valid_o) $display("[TB] Multiple sets: set2_base hit");
        else $display("[TB] ERROR: Multiple sets: set2_base miss");
        pc_i = set3_base; valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
        if (hit_o && valid_o) $display("[TB] Multiple sets: set3_base hit");
        else $display("[TB] ERROR: Multiple sets: set3_base miss");

        // Test 6: Sequential line fills
        $display("[TB] Test 6: Sequential line fills");
        for (int i = 0; i < 4; i++) begin
            pc_i = 32'h4000_0000 + i * LINE_SIZE;
            valid_i = 1; @(posedge clk); valid_i = 0;
            wait (mem_arvalid_o); mem_arready_i = 1; @(posedge clk); mem_arready_i = 0;
            repeat (LINE_SIZE/4) begin mem_rvalid_i = 1; mem_rdata_i = $random; @(posedge clk); end
            mem_rvalid_i = 0; wait (ready_o);
        end
        // Re-access all, should be hits
        for (int i = 0; i < 4; i++) begin
            pc_i = 32'h4000_0000 + i * LINE_SIZE;
            valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
            if (hit_o && valid_o) $display("[TB] Sequential: Hit for addr %h", pc_i);
            else $display("[TB] ERROR: Sequential: Miss for addr %h", pc_i);
        end

        // Test 7: Edge cases (boundary, flush during fill)
        $display("[TB] Test 7: Edge cases");
        // Boundary access
        pc_i = 32'hFFFF_FFE0; // Last line in 32-bit address space
        valid_i = 1; @(posedge clk); valid_i = 0;
        wait (mem_arvalid_o); mem_arready_i = 1; @(posedge clk); mem_arready_i = 0;
        repeat (LINE_SIZE/4) begin mem_rvalid_i = 1; mem_rdata_i = $random; @(posedge clk); end
        mem_rvalid_i = 0; wait (ready_o);
        pc_i = 32'hFFFF_FFE0; valid_i = 1; @(posedge clk); valid_i = 0; @(posedge clk);
        if (hit_o && valid_o) $display("[TB] Edge: Boundary hit");
        else $display("[TB] ERROR: Edge: Boundary miss");
        // Flush during fill
        pc_i = 32'h5000_0000; valid_i = 1; @(posedge clk); valid_i = 0;
        wait (mem_arvalid_o); mem_arready_i = 1; @(posedge clk); mem_arready_i = 0;
        // Start fill, then flush
        mem_rvalid_i = 1; mem_rdata_i = $random; @(posedge clk);
        flush_i = 1; @(posedge clk); flush_i = 0;
        mem_rvalid_i = 0; wait (flush_done_o);
        $display("[TB] Edge: Flushed during fill");
        // Should miss again
        pc_i = 32'h5000_0000; valid_i = 1; @(posedge clk); valid_i = 0;
        wait (mem_arvalid_o); $display("[TB] Edge: Miss after flush during fill as expected");
        mem_arready_i = 1; repeat (LINE_SIZE/4) begin mem_rvalid_i = 1; mem_rdata_i = $random; @(posedge clk); end
        mem_rvalid_i = 0; mem_arready_i = 0; wait (ready_o);
        $display("[TB] Edge: Line refilled after flush during fill");

        // Finish
        $display("[TB] All tests complete");
        $finish;
    end

endmodule : icache_tb

`default_nettype wire 