'module test_wrapper; rtl_core_riscv_core_sv dut(); endmodule' 
