//=============================================================================
// Company: Sondrel Ltd
// Author: DesignAI (designai@sondrel.com)
// Created: 2025-06-27
//
// File: l2_cache.sv
// Module: l2_cache
//
// Project Name: RISC-V RV32IM Core
// Target Devices: ASIC/FPGA
// Verification Status: Not Verified
// Quality Status: Revised Draft
//
// Description:
//   A unified, 8-way set-associative L2 cache for the multi-core system.
//   It serves requests from the L1 caches, maintains coherency via the MESI
//   protocol by interacting with a snooping coherency controller, and
//   forwards misses to the L3 cache. It uses a true LRU replacement policy
//   implemented with a priority encoder based on an internal bit matrix.
//=============================================================================

`timescale 1ns/1ps
`default_nettype none




// AI_TAG: FEATURE - Unified L2 cache for instructions and data.
// AI_TAG: FEATURE - 8-way set-associative with true LRU replacement policy.
// AI_TAG: FEATURE - Maintains MESI coherency across L1 caches.
// AI_TAG: FEATURE - Handles snoop requests from the coherency controller.
// AI_TAG: INTERNAL_BLOCK - RequestArbiter - Round-robin arbiter for L1 requests.
// AI_TAG: INTERNAL_BLOCK - CacheControllerFSM - Main FSM for handling cache requests (hits/misses).
// AI_TAG: INTERNAL_BLOCK - SnoopLogic - Logic to handle incoming snoop requests.
// AI_TAG: INTERNAL_BLOCK - StorageArrays - Tag, Data, and State arrays.
// AI_TAG: INTERNAL_BLOCK - LRU_Logic - Per-set LRU state machine instances.

module l2_cache #(
    parameter integer L2_CACHE_SIZE   = DEFAULT_L2_CACHE_SIZE,     // AI_TAG: PARAM_DESC - L2 cache size in bytes (256KB)
                                                         // AI_TAG: PARAM_USAGE - Determines total cache capacity
                                                         // AI_TAG: PARAM_CONSTRAINTS - Must be power of 2, minimum 64KB
    parameter integer CACHE_LINE_SIZE = DEFAULT_CACHE_LINE_SIZE,             // AI_TAG: PARAM_DESC - Cache line size in bytes (64 Bytes)
                                                         // AI_TAG: PARAM_USAGE - Must match L1 cache line size for coherency
                                                         // AI_TAG: PARAM_CONSTRAINTS - Must be power of 2, typically 32 or 64 bytes
    parameter integer NUM_WAYS        = DEFAULT_L2_NUM_WAYS,              // AI_TAG: PARAM_DESC - Number of ways for set-associativity
                                                         // AI_TAG: PARAM_USAGE - Higher associativity reduces conflict misses
                                                         // AI_TAG: PARAM_CONSTRAINTS - Must be power of 2, typically 4-16
    parameter integer NUM_CORES       = MAX_CORES, // AI_TAG: PARAM_DESC - Number of CPU cores to serve
                                                           // AI_TAG: PARAM_USAGE - Determines interface array sizes
                                                           // AI_TAG: PARAM_CONSTRAINTS - Must match system configuration
    parameter integer DATA_WIDTH      = XLEN,          // AI_TAG: PARAM_DESC - Data bus width
                                                        // AI_TAG: PARAM_USAGE - Must match core data width
                                                        // AI_TAG: PARAM_CONSTRAINTS - Must be XLEN (32 or 64)
    parameter integer ADDR_WIDTH      = ADDR_WIDTH, // AI_TAG: PARAM_DESC - Address bus width
                                                        // AI_TAG: PARAM_USAGE - Determines addressable memory space
                                                        // AI_TAG: PARAM_CONSTRAINTS - Typically 32 or 64 bits
    parameter integer PREFETCH_DEPTH = DEFAULT_L2_PREFETCH_DEPTH,        // How many lines to prefetch ahead
    parameter integer STRIDE_TABLE_SIZE = DEFAULT_L2_STRIDE_TABLE_SIZE,    // Number of stride prediction entries
    parameter integer CONFIDENCE_THRESHOLD = DEFAULT_L2_PREFETCH_CONFIDENCE_THRESHOLD  // Minimum confidence for prefetch
) (
    input  logic clk_i,    // AI_TAG: PORT_DESC - System clock
                           // AI_TAG: PORT_CLK_DOMAIN - clk_i
    input  logic rst_ni,   // AI_TAG: PORT_DESC - Asynchronous active-low reset
                           // AI_TAG: PORT_CLK_DOMAIN - clk_i (async assert)
                           // AI_TAG: PORT_TIMING - Asynchronous

    // Interface to L1 caches (one per core)
    // AI_TAG: IF_TYPE - memory_req_rsp_if (slave)
    // AI_TAG: IF_MODPORT - slave
    // AI_TAG: IF_DESC - Array of interfaces for requests from each L1 cache.
    // AI_TAG: IF_DATA_WIDTHS - Data: DATA_WIDTH, Addr: ADDR_WIDTH
    // AI_TAG: IF_CLOCKING - clk_i
    // AI_TAG: IF_RESET - rst_ni
    memory_req_rsp_if.slave l1_if [NUM_CORES],

    // Interface to L3 cache / Main Memory
    // AI_TAG: IF_TYPE - memory_req_rsp_if (master)
    // AI_TAG: IF_MODPORT - master
    // AI_TAG: IF_DESC - Interface for fetching/writing back data from/to the next memory level.
    // AI_TAG: IF_DATA_WIDTHS - Data: CACHE_LINE_SIZE*8, Addr: ADDR_WIDTH
    // AI_TAG: IF_CLOCKING - clk_i
    // AI_TAG: IF_RESET - rst_ni
    memory_req_rsp_if.master l3_if,

    // Interface to Coherency Controller
    // AI_TAG: IF_TYPE - cache_coherency_if
    // AI_TAG: IF_MODPORT - l2_cache_port
    // AI_TAG: IF_DESC - Interface for snoop requests and coherency management.
    // AI_TAG: IF_CLOCKING - clk_i
    // AI_TAG: IF_RESET - rst_ni
    cache_coherency_if.l2_cache_port coherency_if,

    // Performance Monitoring
    // AI_TAG: PORT_DESC - l1_miss_o - Pulses high for one cycle on an L1 miss for the corresponding core.
    output logic [NUM_CORES-1:0] l1_miss_o
);

    // AI_TAG: CLOCK_SOURCE - clk_i - System clock from clock manager
    // AI_TAG: CLOCK_FREQUENCY_TARGET - clk_i - Up to 1GHz for ASIC, 400MHz for FPGA
    // AI_TAG: RESET_STRATEGY_NOTE - rst_ni is asynchronously asserted and synchronously de-asserted to clk_i
    // AI_TAG: RESET_SYNC_STAGES - rst_ni - 2

    //-----
    // Local Parameters
    //-----
    localparam integer NUM_SETS    = L2_CACHE_SIZE / (CACHE_LINE_SIZE * NUM_WAYS);
    localparam integer OFFSET_BITS = $clog2(CACHE_LINE_SIZE);
    localparam integer INDEX_BITS  = $clog2(NUM_SETS);
    localparam integer TAG_BITS    = ADDR_WIDTH - INDEX_BITS - OFFSET_BITS;
    localparam integer WAY_BITS    = $clog2(NUM_WAYS);
    localparam integer LRU_WIDTH   = (NUM_WAYS * (NUM_WAYS - 1)) / 2;
    localparam integer CORE_ID_BITS = $clog2(NUM_CORES);

    //---------------------------------------------------------------------------
    // L2 Cache Storage Arrays
    //---------------------------------------------------------------------------
    // AI_TAG: INTERNAL_STORAGE - l2_tags_q - Stores the tag for each cache line.
    // AI_TAG: INTERNAL_STORAGE_TYPE - l2_tags_q - SRAM/Register arrays
    // AI_TAG: INTERNAL_STORAGE_ACCESS - l2_tags_q - Read/write by cache controller FSM
    logic [TAG_BITS-1:0]            l2_tags_q  [NUM_SETS-1:0][NUM_WAYS-1:0];
    
    // AI_TAG: INTERNAL_STORAGE - l2_data_q - Stores the actual data for each cache line.
    // AI_TAG: INTERNAL_STORAGE_TYPE - l2_data_q - SRAM arrays
    // AI_TAG: INTERNAL_STORAGE_ACCESS - l2_data_q - Read/write by cache controller FSM
    logic [CACHE_LINE_SIZE*8-1:0]   l2_data_q  [NUM_SETS-1:0][NUM_WAYS-1:0];
    
    // AI_TAG: INTERNAL_STORAGE - l2_state_q - Stores the MESI state for each cache line.
    // AI_TAG: INTERNAL_STORAGE_TYPE - l2_state_q - Register arrays
    // AI_TAG: INTERNAL_STORAGE_ACCESS - l2_state_q - Read/write by coherency and cache logic
    cache_state_t                   l2_state_q [NUM_SETS-1:0][NUM_WAYS-1:0];
    
    // AI_TAG: INTERNAL_STORAGE - l2_lru_q - Stores the LRU state for each set.
    // AI_TAG: INTERNAL_STORAGE_TYPE - l2_lru_q - Register arrays
    // AI_TAG: INTERNAL_STORAGE_ACCESS - l2_lru_q - Read/write by LRU management logic
    logic [LRU_WIDTH-1:0]           l2_lru_q   [NUM_SETS-1:0];
    logic [LRU_WIDTH-1:0]           l2_lru_ns;

    //---------------------------------------------------------------------------
    // FSM for Cache Controller Logic
    //---------------------------------------------------------------------------
    // AI_TAG: FSM_NAME - cache_controller_fsm
    // AI_TAG: FSM_PURPOSE - cache_controller_fsm - Controls cache operations for hits, misses, and coherency
    // AI_TAG: FSM_ENCODING - cache_controller_fsm - one-hot for performance
    // AI_TAG: FSM_RESET_STATE - cache_controller_fsm - IDLE
    // AI_TAG: FSM_INPUT_CONDITIONS - cache_controller_fsm - l1_req_valid, l3_rsp_valid, snoop_req
    typedef enum logic [3:0] {
        IDLE            = 4'b0001,  // AI_TAG: FSM_STATE - IDLE - Waiting for L1 requests
        TAG_CHECK       = 4'b0010,  // AI_TAG: FSM_STATE - TAG_CHECK - Checking tags for hit/miss
        READ_HIT        = 4'b0100,  // AI_TAG: FSM_STATE - READ_HIT - Servicing read hit
        WRITE_HIT       = 4'b1000,  // AI_TAG: FSM_STATE - WRITE_HIT - Servicing write hit
        EVICT_WRITEBACK = 4'b0011,  // AI_TAG: FSM_STATE - EVICT_WRITEBACK - Writing back dirty victim
        FETCH_L3        = 4'b0101,  // AI_TAG: FSM_STATE - FETCH_L3 - Fetching missing line from L3
        REFILL_L2       = 4'b1001,  // AI_TAG: FSM_STATE - REFILL_L2 - Installing fetched line
        RESPOND         = 4'b0110   // AI_TAG: FSM_STATE - RESPOND - Sending response to L1
    } cache_state_e;

    cache_state_e current_state_r, next_state_c;

    // AI_TAG: INTERNAL_LOGIC - Miss tracking for performance monitoring
    logic [NUM_CORES-1:0] l1_miss_w;

    // AI_TAG: FSM_OUTPUT_ACTIONS - cache_controller_fsm - IDLE - All interfaces idle, ready for new requests
    // AI_TAG: FSM_OUTPUT_ACTIONS - cache_controller_fsm - TAG_CHECK - Tag comparison active, way selection logic enabled
    // AI_TAG: FSM_OUTPUT_ACTIONS - cache_controller_fsm - READ_HIT - Data output enabled, LRU update triggered
    // AI_TAG: FSM_OUTPUT_ACTIONS - cache_controller_fsm - WRITE_HIT - Data write enabled, state update to Modified
    // AI_TAG: FSM_OUTPUT_ACTIONS - cache_controller_fsm - EVICT_WRITEBACK - L3 write request active with victim data
    // AI_TAG: FSM_OUTPUT_ACTIONS - cache_controller_fsm - FETCH_L3 - L3 read request active for missing line
    // AI_TAG: FSM_OUTPUT_ACTIONS - cache_controller_fsm - REFILL_L2 - Cache arrays write enabled, LRU update
    // AI_TAG: FSM_OUTPUT_ACTIONS - cache_controller_fsm - RESPOND - L1 response valid with result data

    // Registers for active request
    memory_req_t      active_req_r;
    logic [CORE_ID_BITS-1:0] active_core_id_r;
    logic [WAY_BITS-1:0]     hit_way_r;
    logic             is_hit_r;
    logic [WAY_BITS-1:0]     victim_way_r;
    logic [CACHE_LINE_SIZE*8-1:0] victim_data_r;
    logic [ADDR_WIDTH-1:0]        victim_addr_r;

    // Address decoding
    logic [INDEX_BITS-1:0] index_c;
    logic [TAG_BITS-1:0]   tag_c;
    logic [OFFSET_BITS-1:0] offset_c;

    assign index_c  = active_req_r.addr[OFFSET_BITS +: INDEX_BITS];
    assign tag_c    = active_req_r.addr[ADDR_WIDTH-1 -: TAG_BITS];
    assign offset_c = active_req_r.addr[OFFSET_BITS-1:0];

    //---------------------------------------------------------------------------
    // Hardware Cache Prefetcher - Next-Line and Stride Prediction
    //---------------------------------------------------------------------------
    // AI_TAG: PERFORMANCE_FEATURE - Hardware prefetcher for improved cache performance
    // AI_TAG: FEATURE - Next-line prefetching and stride-based prediction
    
    // Prefetcher Configuration
    localparam integer PREFETCH_DEPTH = DEFAULT_L2_PREFETCH_DEPTH;        // How many lines to prefetch ahead
    localparam integer STRIDE_TABLE_SIZE = DEFAULT_L2_STRIDE_TABLE_SIZE;    // Number of stride prediction entries
    localparam integer CONFIDENCE_THRESHOLD = DEFAULT_L2_PREFETCH_CONFIDENCE_THRESHOLD;  // Minimum confidence for prefetch
    
    // Stride Prediction Table Entry
    typedef struct packed {
        logic [ADDR_WIDTH-1:0] last_addr;
        logic [ADDR_WIDTH-1:0] stride;
        logic [2:0] confidence;
        logic [CORE_ID_BITS-1:0] core_id;
        logic valid;
    } stride_entry_t;
    
    stride_entry_t stride_table [STRIDE_TABLE_SIZE-1:0];
    logic [$clog2(STRIDE_TABLE_SIZE)-1:0] stride_table_ptr_r;
    
    // Prefetch Request Generation
    logic prefetch_req_valid_c;
    logic [ADDR_WIDTH-1:0] prefetch_addr_c;
    logic [CORE_ID_BITS-1:0] prefetch_core_c;
    logic prefetch_granted_r;
    
    // Prefetch FSM
    typedef enum logic [1:0] {
        PREFETCH_IDLE     = 2'b00,
        PREFETCH_GENERATE = 2'b01,
        PREFETCH_ISSUE    = 2'b10,
        PREFETCH_WAIT     = 2'b11
    } prefetch_state_e;
    
    prefetch_state_e prefetch_state_r;
    
    //-----
    // Stride Prediction and Prefetch Generation
    //-----
    always_ff @(posedge clk_i or negedge rst_ni) begin : proc_prefetcher
        if (!rst_ni) begin
            for (int i = 0; i < STRIDE_TABLE_SIZE; i++) begin
                stride_table[i] <= '0;
            end
            stride_table_ptr_r <= '0;
            prefetch_state_r <= PREFETCH_IDLE;
            prefetch_granted_r <= 1'b0;
        end else begin
            // Update stride prediction table on L1 requests
            if (current_state_r == TAG_CHECK && is_hit_r) begin
                logic [$clog2(STRIDE_TABLE_SIZE)-1:0] match_idx;
                logic match_found = 1'b0;
                
                // Look for existing entry for this core
                for (int i = 0; i < STRIDE_TABLE_SIZE; i++) begin
                    if (stride_table[i].valid && 
                        stride_table[i].core_id == active_core_id_r && 
                        !match_found) begin
                        match_idx = i;
                        match_found = 1'b1;
                    end
                end
                
                if (match_found) begin
                    // Update existing entry
                    logic [ADDR_WIDTH-1:0] new_stride = active_req_r.addr - stride_table[match_idx].last_addr;
                    
                    if (new_stride == stride_table[match_idx].stride) begin
                        // Stride confirmed, increase confidence
                        if (stride_table[match_idx].confidence < 7) begin
                            stride_table[match_idx].confidence <= stride_table[match_idx].confidence + 1;
                        end
                    end else begin
                        // New stride pattern
                        stride_table[match_idx].stride <= new_stride;
                        stride_table[match_idx].confidence <= 1;
                    end
                    stride_table[match_idx].last_addr <= active_req_r.addr;
                end else begin
                    // Create new entry
                    stride_table[stride_table_ptr_r] <= '{
                        last_addr: active_req_r.addr,
                        stride: CACHE_LINE_SIZE, // Default to next-line
                        confidence: 1,
                        core_id: active_core_id_r,
                        valid: 1'b1
                    };
                    stride_table_ptr_r <= stride_table_ptr_r + 1;
                end
            end
            
            // Prefetch State Machine
            case (prefetch_state_r)
                PREFETCH_IDLE: begin
                    prefetch_granted_r <= 1'b0;
                    // Trigger prefetch on cache miss
                    if (current_state_r == FETCH_L3 && l3_if.req_ready) begin
                        prefetch_state_r <= PREFETCH_GENERATE;
                    end
                end
                
                PREFETCH_GENERATE: begin
                    // Check if we should prefetch
                    prefetch_state_r <= PREFETCH_ISSUE;
                end
                
                PREFETCH_ISSUE: begin
                    // Issue prefetch request if L3 is ready and no higher priority traffic
                    if (l3_if.req_ready && current_state_r == IDLE) begin
                        prefetch_granted_r <= 1'b1;
                        prefetch_state_r <= PREFETCH_WAIT;
                    end
                end
                
                PREFETCH_WAIT: begin
                    // Wait for prefetch completion
                    if (l3_if.rsp_valid && prefetch_granted_r) begin
                        prefetch_granted_r <= 1'b0;
                        prefetch_state_r <= PREFETCH_IDLE;
                    end
                end
            endcase
        end
    end
    
    //-----
    // Prefetch Address Generation
    //-----
    always_comb begin : proc_prefetch_addr_gen
        prefetch_req_valid_c = 1'b0;
        prefetch_addr_c = '0;
        prefetch_core_c = '0;
        
        if (prefetch_state_r == PREFETCH_ISSUE) begin
            // Find highest confidence stride entry
            logic [2:0] best_confidence = '0;
            logic [$clog2(STRIDE_TABLE_SIZE)-1:0] best_idx = '0;
            logic prefetch_candidate_found = 1'b0;
            
            for (int i = 0; i < STRIDE_TABLE_SIZE; i++) begin
                if (stride_table[i].valid && 
                    stride_table[i].confidence >= CONFIDENCE_THRESHOLD &&
                    stride_table[i].confidence > best_confidence) begin
                    best_confidence = stride_table[i].confidence;
                    best_idx = i;
                    prefetch_candidate_found = 1'b1;
                end
            end
            
            if (prefetch_candidate_found) begin
                prefetch_req_valid_c = 1'b1;
                prefetch_addr_c = stride_table[best_idx].last_addr + stride_table[best_idx].stride;
                prefetch_core_c = stride_table[best_idx].core_id;
            end
        end
    end

    // LRU management signals
    logic [WAY_BITS-1:0]  lru_victim_way_c;
    logic                 lru_update_en_c;
    logic [WAY_BITS-1:0]  lru_update_way_c;

    // Round-robin arbiter for L1 requests
    logic [CORE_ID_BITS-1:0] arbiter_grant_r;
    logic                    arbiter_grant_valid_c;

    //---------------------------------------------------------------------------
    // Round-Robin Arbiter for L1 Requests
    //---------------------------------------------------------------------------
    always_ff @(posedge clk_i or negedge rst_ni) begin : proc_arbiter
        if (!rst_ni) begin
            arbiter_grant_r <= '0;
        end else if (current_state_r == IDLE && arbiter_grant_valid_c) begin
            arbiter_grant_r <= arbiter_grant_r + 1;
        end
    end

    always_comb begin : proc_arbiter_logic
        arbiter_grant_valid_c = 1'b0;
        
        // Find next requesting core starting from current grant pointer
        for (int i = 0; i < NUM_CORES; i++) begin
            logic [CORE_ID_BITS-1:0] core_idx = (arbiter_grant_r + i) % NUM_CORES;
            if (l1_if[core_idx].req_valid) begin
                arbiter_grant_valid_c = 1'b1;
                break;
            end
        end
    end

    //---------------------------------------------------------------------------
    // LRU Management Logic
    //---------------------------------------------------------------------------
    genvar i;
    generate
        for (i = 0; i < NUM_SETS; i++) begin : gen_lru
            matrix_lru #(
                .NUM_WAYS(NUM_WAYS)
            ) u_matrix_lru (
                .clk_i        (clk_i),
                .rst_ni       (rst_ni),
                .update_en_i  (lru_update_en_c && (index_c == i)),
                .update_way_i (lru_update_way_c),
                .lru_way_o    (lru_victim_way_c),
                .lru_state_i  (l2_lru_q[i]),
                .lru_state_o  (l2_lru_ns)
            );
        end
    endgenerate

    //---------------------------------------------------------------------------
    // Main Cache Controller FSM
    //---------------------------------------------------------------------------
    // AI_TAG: FSM_TRANSITION - cache_controller_fsm: IDLE -> TAG_CHECK when (arbiter_grant_valid_c)
    // AI_TAG: FSM_TRANSITION - cache_controller_fsm: TAG_CHECK -> READ_HIT when (is_hit_r && !active_req_r.write)
    // AI_TAG: FSM_TRANSITION - cache_controller_fsm: TAG_CHECK -> WRITE_HIT when (is_hit_r && active_req_r.write)
    // AI_TAG: FSM_TRANSITION - cache_controller_fsm: TAG_CHECK -> EVICT_WRITEBACK when (!is_hit_r && victim_needs_writeback)
    // AI_TAG: FSM_TRANSITION - cache_controller_fsm: TAG_CHECK -> FETCH_L3 when (!is_hit_r && !victim_needs_writeback)
    // AI_TAG: FSM_TRANSITION - cache_controller_fsm: EVICT_WRITEBACK -> FETCH_L3 when (l3_if.req_ready)
    // AI_TAG: FSM_TRANSITION - cache_controller_fsm: FETCH_L3 -> REFILL_L2 when (l3_if.req_ready)
    // AI_TAG: FSM_TRANSITION - cache_controller_fsm: REFILL_L2 -> RESPOND when (l3_if.rsp_valid)
    // AI_TAG: FSM_TRANSITION - cache_controller_fsm: RESPOND -> IDLE when (l1_response_accepted)

    always_ff @(posedge clk_i or negedge rst_ni) begin : proc_cache_fsm_reg
        if (!rst_ni) begin
            current_state_r <= IDLE;
            // Reset all cache arrays
            for (int i = 0; i < NUM_SETS; i++) begin
                for (int j = 0; j < NUM_WAYS; j++) begin
                    l2_tags_q[i][j] <= '0;
                    l2_data_q[i][j] <= '0;
                    l2_state_q[i][j] <= CACHE_INVALID; // Invalid state
                end
                l2_lru_q[i] <= '0;
            end
            // Reset FSM registers
            active_req_r <= '0;
            active_core_id_r <= '0;
            hit_way_r <= '0;
            is_hit_r <= '0;
            victim_way_r <= '0;
            victim_data_r <= '0;
            victim_addr_r <= '0;
        end else begin
            current_state_r <= next_state_c;
            
            // Update LRU when enabled
            if (lru_update_en_c) begin
                l2_lru_q[index_c] <= l2_lru_ns;
            end
            
            // Register active request when transitioning from IDLE
            if (current_state_r == IDLE && next_state_c == TAG_CHECK) begin
                logic [CORE_ID_BITS-1:0] granted_core = (arbiter_grant_r + 0) % NUM_CORES;
                for (int k = 0; k < NUM_CORES; k++) begin
                    logic [CORE_ID_BITS-1:0] core_idx = (arbiter_grant_r + k) % NUM_CORES;
                    if (l1_if[core_idx].req_valid) begin
                        granted_core = core_idx;
                        break;
                    end
                end
                active_req_r <= l1_if[granted_core].req;
                active_core_id_r <= granted_core;
            end
            
            // Update cache arrays during refill
            if (current_state_r == REFILL_L2 && l3_if.rsp_valid) begin
                l2_tags_q[index_c][victim_way_r] <= tag_c;
                l2_data_q[index_c][victim_way_r] <= l3_if.rsp.data;
                l2_state_q[index_c][victim_way_r] <= active_req_r.write ? CACHE_MODIFIED : CACHE_SHARED;
            end
            
            // Update cache state during write hit
            if (current_state_r == WRITE_HIT) begin
                l2_state_q[index_c][hit_way_r] <= CACHE_MODIFIED;
                // Update specific bytes in cache line
                for (int byte_idx = 0; byte_idx < DATA_WIDTH/8; byte_idx++) begin
                    if (active_req_r.strb[byte_idx]) begin
                        l2_data_q[index_c][hit_way_r][offset_c*8 + byte_idx*8 +: 8] <= 
                            active_req_r.data[byte_idx*8 +: 8];
                    end
                end
            end
        end
    end

    always_comb begin : proc_cache_fsm_logic
        next_state_c = current_state_r;
        
        // Default output assignments
        for(int j=0; j<NUM_CORES; j++) begin
            l1_if[j].req_ready = 1'b0;
            l1_if[j].rsp_valid = 1'b0;
            l1_if[j].rsp = '0;
        end
        l3_if.req_valid = 1'b0;
        l3_if.req = '0;
        l3_if.rsp_ready = 1'b1; // Always ready to accept L3 responses

        lru_update_en_c = 1'b0;
        lru_update_way_c = '0;
        l1_miss_w = '0;

        case (current_state_r)
            IDLE: begin
                if (arbiter_grant_valid_c) begin
                    // Accept request from granted core
                    logic [CORE_ID_BITS-1:0] granted_core = (arbiter_grant_r + 0) % NUM_CORES;
                    for (int k = 0; k < NUM_CORES; k++) begin
                        logic [CORE_ID_BITS-1:0] core_idx = (arbiter_grant_r + k) % NUM_CORES;
                        if (l1_if[core_idx].req_valid) begin
                            granted_core = core_idx;
                            break;
                        end
                    end
                    l1_if[granted_core].req_ready = 1'b1;
                    next_state_c = TAG_CHECK;
                end else if (prefetch_req_valid_c && l3_if.req_ready) begin
                    // Handle prefetch request when no other traffic
                    l3_if.req_valid = 1'b1;
                    l3_if.req.addr = {prefetch_addr_c[ADDR_WIDTH-1:OFFSET_BITS], {OFFSET_BITS{1'b0}}};
                    l3_if.req.data = '0;
                    l3_if.req.write = 1'b0;
                    l3_if.req.strb = '1;
                    l3_if.req.id = 8'hFF; // Special prefetch ID
                    l3_if.req.last = 1'b1;
                    // Stay in IDLE for prefetch - no state change needed
                end
            end

            TAG_CHECK: begin
                logic has_invalid_way_c;
                logic [WAY_BITS-1:0] invalid_way_idx_c;
                
                is_hit_r = 1'b0;
                has_invalid_way_c = 1'b0;
                invalid_way_idx_c = '0;

                // Check for hit and find invalid way
                for (int j = 0; j < NUM_WAYS; j++) begin
                    if (l2_state_q[index_c][j] == CACHE_INVALID) begin
                        if (!has_invalid_way_c) begin // Take first invalid way found
                            has_invalid_way_c = 1'b1;
                            invalid_way_idx_c = WAY_BITS'(j);
                        end
                    end else if (l2_tags_q[index_c][j] == tag_c) begin
                        is_hit_r = 1'b1;
                        hit_way_r = WAY_BITS'(j);
                    end
                end
                
                if (is_hit_r) begin
                    // Cache hit - update LRU and proceed based on operation
                    lru_update_en_c = 1'b1;
                    lru_update_way_c = hit_way_r;
                    next_state_c = active_req_r.write ? WRITE_HIT : READ_HIT;
                end else begin
                    // Cache miss - determine victim and check if writeback needed
                    victim_way_r = has_invalid_way_c ? invalid_way_idx_c : lru_victim_way_c;
                    l1_miss_w[active_core_id_r] = 1'b1; // Signal miss for this core
                    
                    if (l2_state_q[index_c][victim_way_r] == CACHE_MODIFIED && !has_invalid_way_c) begin
                        // Victim is dirty and needs writeback
                        victim_data_r = l2_data_q[index_c][victim_way_r];
                        victim_addr_r = {l2_tags_q[index_c][victim_way_r], index_c, {OFFSET_BITS{1'b0}}};
                        next_state_c = EVICT_WRITEBACK;
                    end else begin
                        // No writeback needed, go directly to fetch
                        next_state_c = FETCH_L3;
                    end
                end
            end

            READ_HIT: begin
                next_state_c = RESPOND;
            end
            
            WRITE_HIT: begin
                next_state_c = RESPOND;
            end

            EVICT_WRITEBACK: begin
                // Setup L3 write request for victim line
                l3_if.req_valid = 1'b1;
                l3_if.req.addr = victim_addr_r;
                l3_if.req.data = victim_data_r;
                l3_if.req.write = 1'b1;
                l3_if.req.strb = '1; // Write entire cache line
                l3_if.req.id = active_req_r.id;
                l3_if.req.last = 1'b1;
                
                if (l3_if.req_ready) begin
                    next_state_c = FETCH_L3;
                end
            end

            FETCH_L3: begin
                // Setup L3 read request for missing line
                l3_if.req_valid = 1'b1;
                l3_if.req.addr = {tag_c, index_c, {OFFSET_BITS{1'b0}}}; // Aligned address
                l3_if.req.data = '0;
                l3_if.req.write = 1'b0;
                l3_if.req.strb = '1; // Read entire cache line
                l3_if.req.id = active_req_r.id;
                l3_if.req.last = 1'b1;
                
                if (l3_if.req_ready) begin
                    next_state_c = REFILL_L2;
                end
            end

            REFILL_L2: begin
                if (l3_if.rsp_valid) begin
                    // Cache line will be updated in sequential block
                    lru_update_en_c = 1'b1;
                    lru_update_way_c = victim_way_r;
                    next_state_c = RESPOND;
                end
            end
            
            RESPOND: begin
                // Send response to requesting L1 cache
                l1_if[active_core_id_r].rsp_valid = 1'b1;
                l1_if[active_core_id_r].rsp.id = active_req_r.id;
                l1_if[active_core_id_r].rsp.error = 1'b0;
                l1_if[active_core_id_r].rsp.last = 1'b1;
                
                if (active_req_r.write) begin
                    // Write response - no data
                    l1_if[active_core_id_r].rsp.data = '0;
                end else begin
                    // Read response - extract requested data from cache line
                    if (current_state_r == READ_HIT) begin
                        // Extract data from hit way
                        l1_if[active_core_id_r].rsp.data = 
                            l2_data_q[index_c][hit_way_r][offset_c*8 +: DATA_WIDTH];
                    end else begin
                        // Extract data from refilled line
                        l1_if[active_core_id_r].rsp.data = 
                            l3_if.rsp.data[offset_c*8 +: DATA_WIDTH];
                    end
                end
                
                if (l1_if[active_core_id_r].rsp_ready) begin
                    next_state_c = IDLE;
                end
            end

            default: begin
                next_state_c = IDLE;
            end
        endcase
    end
    
    // Register the miss signal to create a single-cycle pulse
    logic [NUM_CORES-1:0] l1_miss_r;
    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            l1_miss_r <= '0;
        end else begin
            l1_miss_r <= l1_miss_w;
        end
    end
    assign l1_miss_o = l1_miss_r;

    //------------------------------------------------------------------------- 
    // Snoop Handling Logic for Cache Coherency
    //-------------------------------------------------------------------------
    // AI_TAG: SNOOP_HANDLER - Handles coherency snoops from other caches
    // AI_TAG: FEATURE - MESI protocol snoop response handling
    always_ff @(posedge clk_i or negedge rst_ni) begin : proc_snoop_handler
        if (!rst_ni) begin
            // Reset snoop response signals
            for (int i = 0; i < NUM_CORES; i++) begin
                coherency_if.snoop_rsp_valid[i] <= 1'b0;
                coherency_if.snoop_rsp_data_valid[i] <= 1'b0;
                coherency_if.snoop_rsp_data[i] <= '0;
            end
        end else begin
            // Handle snoop requests from cache coherency controller
            for (int i = 0; i < NUM_CORES; i++) begin
                if (coherency_if.snoop_valid[i]) begin
                    logic [INDEX_BITS-1:0] snoop_index = 
                        coherency_if.snoop_addr[i][OFFSET_BITS +: INDEX_BITS];
                    logic [TAG_BITS-1:0] snoop_tag = 
                        coherency_if.snoop_addr[i][ADDR_WIDTH-1 -: TAG_BITS];
                    logic snoop_hit = 1'b0;
                    logic [WAY_BITS-1:0] snoop_way = '0;
                    
                    // Check for hit in all ways
                    for (int j = 0; j < NUM_WAYS; j++) begin
                        if (l2_tags_q[snoop_index][j] == snoop_tag && 
                            l2_state_q[snoop_index][j] != CACHE_INVALID) begin
                            snoop_hit = 1'b1;
                            snoop_way = WAY_BITS'(j);
                            break;
                        end
                    end
                    
                    // Process snoop based on type
                    case (coherency_if.snoop_type[i])
                        COHERENCY_REQ_INVALIDATE: begin
                            if (snoop_hit) begin
                                l2_state_q[snoop_index][snoop_way] <= CACHE_INVALID;
                            end
                            coherency_if.snoop_rsp_valid[i] <= 1'b1;
                            coherency_if.snoop_rsp_data_valid[i] <= 1'b0;
                        end
                        
                        COHERENCY_REQ_READ: begin
                            if (snoop_hit) begin
                                coherency_if.snoop_rsp_data[i] <= l2_data_q[snoop_index][snoop_way];
                                coherency_if.snoop_rsp_data_valid[i] <= 1'b1;
                                // Downgrade state if in Modified
                                if (l2_state_q[snoop_index][snoop_way] == CACHE_MODIFIED) begin
                                    l2_state_q[snoop_index][snoop_way] <= CACHE_SHARED;
                                end
                            end else begin
                                coherency_if.snoop_rsp_data_valid[i] <= 1'b0;
                            end
                            coherency_if.snoop_rsp_valid[i] <= 1'b1;
                        end
                        
                        default: begin
                            coherency_if.snoop_rsp_valid[i] <= 1'b1;
                            coherency_if.snoop_rsp_data_valid[i] <= 1'b0;
                        end
                    endcase
                end else begin
                    // Clear response when no snoop
                    coherency_if.snoop_rsp_valid[i] <= 1'b0;
                    coherency_if.snoop_rsp_data_valid[i] <= 1'b0;
                end
            end
        end
    end

    // AI_TAG: ASSERTION - a_cache_hit_exclusive: Cache hit should occur in at most one way
    // AI_TAG: ASSERTION_TYPE - Simulation
    // AI_TAG: ASSERTION_SEVERITY - Error
`ifdef SIMULATION
    always_comb begin : proc_assertions
        // Check that at most one way has a hit for any given address
        if (current_state_r == TAG_CHECK) begin
            logic [NUM_WAYS-1:0] hit_vector;
            for (int j = 0; j < NUM_WAYS; j++) begin
                hit_vector[j] = (l2_tags_q[index_c][j] == tag_c) && 
                               (l2_state_q[index_c][j] != CACHE_INVALID);
            end
            assert ($onehot0(hit_vector)) 
                else $error("Multiple cache ways hit for address %h", active_req_r.addr);
        end
    end
`endif

endmodule : l2_cache

//=============================================================================
// Dependencies:
//   - rtl/core/riscv_config_pkg.sv
//   - rtl/core/riscv_types_pkg.sv
//   - rtl/core/riscv_cache_types_pkg.sv
//   - rtl/core/riscv_mem_types_pkg.sv
//   - rtl/memory/memory_req_rsp_if.sv
//   - rtl/interfaces/cache_coherency_if.sv
//   - rtl/memory/matrix_lru.sv
// Instantiated In:
//   - rtl/core/riscv_core.sv
//   - rtl/memory/controllers/cache_cluster_manager.sv
//   - tb/integration/memory_subsystem_integration_tb.sv
//
// Performance:
//   - Critical Path: Tag comparison and way selection logic
//   - Max Frequency: Target 1GHz ASIC, 400MHz FPGA
//   - Area: ~50K gates for 256KB cache with LRU
//
// Verification Coverage:
//   - Code Coverage: TBD
//   - Functional Coverage: All MESI state transitions
//   - Branch Coverage: All FSM paths and cache scenarios
//
// Synthesis:
//   - Target Technology: ASIC/FPGA
//   - Synthesis Tool: Design Compiler/Quartus
//   - Clock Domains: 1 (clk_i)
//   - Constraints File: l2_cache.sdc
//
// Testing:
//   - Testbench: l2_cache_tb.sv (to be created)
//   - Test Vectors: Multi-core coherency scenarios
//
//----
// Revision History:
// Version | Date       | Author             | Description
//=============================================================================
// 2.0.0   | 2025-01-27 | DesignAI           | Fixed critical issues: syntax errors, completed FSM logic, added proper data handling
// 1.0.0   | 2025-06-28 | DesignAI           | Initial fleshed-out implementation.
// 0.1.0   | 2025-06-27 | DesignAI           | Initial skeleton release
//=============================================================================

`default_nettype wire